--------------------------------------------------------------------------------
--  UMass , Physics Department
--  Guillermo Loustau de Linares
--  gloustau@cern.ch
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger 
--  Module: slc vector processor slope calculator
--  Description:
--
--------------------------------------------------------------------------------
--  Revisions:
--      
--------------------------------------------------------------------------------
library ieee, shared_lib;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;
use shared_lib.config_pkg.all;
 
-- library ucm_lib;
-- use ucm_lib.ucm_pkg.all;
-- use ucm_lib.roi_atan.all;

entity ucm_cvp_atan is
  port (
    clk                 : in std_logic;
    rst                 : in std_logic;
    glob_en             : in std_logic
    
  );
end entity ucm_cvp_atan;

architecture beh of ucm_cvp_atan is
  
begin
  
  
  
end architecture beh;