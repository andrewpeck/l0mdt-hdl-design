--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: slope to angle (mrad) 
--  Multiplier: 100000 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library heg_roi_lib;
use heg_roi_lib.roi_types_pkg.all;

package roi_atan is

  -- add length of constant array
  constant ROM_ATAN_MAX_SIZE : integer := 111638;

  type roi_atan_lut_t is array (integer range <> ) of integer;

  constant ROI_ATAN_MEM : roi_atan_lut_t(0 to ROM_ATAN_MAX_SIZE - 1) := (

        0 to    49 =>    0,
       50 to   149 =>    1,
      150 to   249 =>    2,
      250 to   349 =>    3,
      350 to   449 =>    4,
      450 to   549 =>    5,
      550 to   649 =>    6,
      650 to   749 =>    7,
      750 to   849 =>    8,
      850 to   949 =>    9,
      950 to  1049 =>   10,
     1050 to  1149 =>   11,
     1150 to  1249 =>   12,
     1250 to  1349 =>   13,
     1350 to  1449 =>   14,
     1450 to  1549 =>   15,
     1550 to  1649 =>   16,
     1650 to  1749 =>   17,
     1750 to  1849 =>   18,
     1850 to  1949 =>   19,
     1950 to  2049 =>   20,
     2050 to  2149 =>   21,
     2150 to  2249 =>   22,
     2250 to  2349 =>   23,
     2350 to  2449 =>   24,
     2450 to  2548 =>   25,
     2549 to  2648 =>   26,
     2649 to  2748 =>   27,
     2749 to  2848 =>   28,
     2849 to  2948 =>   29,
     2949 to  3048 =>   30,
     3049 to  3148 =>   31,
     3149 to  3248 =>   32,
     3249 to  3348 =>   33,
     3349 to  3448 =>   34,
     3449 to  3548 =>   35,
     3549 to  3647 =>   36,
     3648 to  3747 =>   37,
     3748 to  3847 =>   38,
     3848 to  3947 =>   39,
     3948 to  4047 =>   40,
     4048 to  4147 =>   41,
     4148 to  4246 =>   42,
     4247 to  4346 =>   43,
     4347 to  4446 =>   44,
     4447 to  4546 =>   45,
     4547 to  4646 =>   46,
     4647 to  4745 =>   47,
     4746 to  4845 =>   48,
     4846 to  4945 =>   49,
     4946 to  5045 =>   50,
     5046 to  5144 =>   51,
     5145 to  5244 =>   52,
     5245 to  5344 =>   53,
     5345 to  5444 =>   54,
     5445 to  5543 =>   55,
     5544 to  5643 =>   56,
     5644 to  5743 =>   57,
     5744 to  5842 =>   58,
     5843 to  5942 =>   59,
     5943 to  6042 =>   60,
     6043 to  6141 =>   61,
     6142 to  6241 =>   62,
     6242 to  6340 =>   63,
     6341 to  6440 =>   64,
     6441 to  6540 =>   65,
     6541 to  6639 =>   66,
     6640 to  6739 =>   67,
     6740 to  6838 =>   68,
     6839 to  6938 =>   69,
     6939 to  7037 =>   70,
     7038 to  7137 =>   71,
     7138 to  7236 =>   72,
     7237 to  7336 =>   73,
     7337 to  7435 =>   74,
     7436 to  7535 =>   75,
     7536 to  7634 =>   76,
     7635 to  7734 =>   77,
     7735 to  7833 =>   78,
     7834 to  7932 =>   79,
     7933 to  8032 =>   80,
     8033 to  8131 =>   81,
     8132 to  8230 =>   82,
     8231 to  8330 =>   83,
     8331 to  8429 =>   84,
     8430 to  8528 =>   85,
     8529 to  8628 =>   86,
     8629 to  8727 =>   87,
     8728 to  8826 =>   88,
     8827 to  8925 =>   89,
     8926 to  9024 =>   90,
     9025 to  9124 =>   91,
     9125 to  9223 =>   92,
     9224 to  9322 =>   93,
     9323 to  9421 =>   94,
     9422 to  9520 =>   95,
     9521 to  9619 =>   96,
     9620 to  9718 =>   97,
     9719 to  9817 =>   98,
     9818 to  9916 =>   99,
     9917 to 10015 =>  100,
    10016 to 10114 =>  101,
    10115 to 10213 =>  102,
    10214 to 10312 =>  103,
    10313 to 10411 =>  104,
    10412 to 10510 =>  105,
    10511 to 10609 =>  106,
    10610 to 10708 =>  107,
    10709 to 10807 =>  108,
    10808 to 10906 =>  109,
    10907 to 11004 =>  110,
    11005 to 11103 =>  111,
    11104 to 11202 =>  112,
    11203 to 11301 =>  113,
    11302 to 11399 =>  114,
    11400 to 11498 =>  115,
    11499 to 11597 =>  116,
    11598 to 11695 =>  117,
    11696 to 11794 =>  118,
    11795 to 11893 =>  119,
    11894 to 11991 =>  120,
    11992 to 12090 =>  121,
    12091 to 12188 =>  122,
    12189 to 12287 =>  123,
    12288 to 12385 =>  124,
    12386 to 12484 =>  125,
    12485 to 12582 =>  126,
    12583 to 12681 =>  127,
    12682 to 12779 =>  128,
    12780 to 12877 =>  129,
    12878 to 12976 =>  130,
    12977 to 13074 =>  131,
    13075 to 13172 =>  132,
    13173 to 13271 =>  133,
    13272 to 13369 =>  134,
    13370 to 13467 =>  135,
    13468 to 13565 =>  136,
    13566 to 13663 =>  137,
    13664 to 13761 =>  138,
    13762 to 13860 =>  139,
    13861 to 13958 =>  140,
    13959 to 14056 =>  141,
    14057 to 14154 =>  142,
    14155 to 14252 =>  143,
    14253 to 14350 =>  144,
    14351 to 14448 =>  145,
    14449 to 14546 =>  146,
    14547 to 14643 =>  147,
    14644 to 14741 =>  148,
    14742 to 14839 =>  149,
    14840 to 14937 =>  150,
    14938 to 15035 =>  151,
    15036 to 15132 =>  152,
    15133 to 15230 =>  153,
    15231 to 15328 =>  154,
    15329 to 15425 =>  155,
    15426 to 15523 =>  156,
    15524 to 15621 =>  157,
    15622 to 15718 =>  158,
    15719 to 15816 =>  159,
    15817 to 15913 =>  160,
    15914 to 16011 =>  161,
    16012 to 16108 =>  162,
    16109 to 16206 =>  163,
    16207 to 16303 =>  164,
    16304 to 16400 =>  165,
    16401 to 16498 =>  166,
    16499 to 16595 =>  167,
    16596 to 16692 =>  168,
    16693 to 16789 =>  169,
    16790 to 16887 =>  170,
    16888 to 16984 =>  171,
    16985 to 17081 =>  172,
    17082 to 17178 =>  173,
    17179 to 17275 =>  174,
    17276 to 17372 =>  175,
    17373 to 17469 =>  176,
    17470 to 17566 =>  177,
    17567 to 17663 =>  178,
    17664 to 17760 =>  179,
    17761 to 17857 =>  180,
    17858 to 17954 =>  181,
    17955 to 18050 =>  182,
    18051 to 18147 =>  183,
    18148 to 18244 =>  184,
    18245 to 18341 =>  185,
    18342 to 18437 =>  186,
    18438 to 18534 =>  187,
    18535 to 18630 =>  188,
    18631 to 18727 =>  189,
    18728 to 18823 =>  190,
    18824 to 18920 =>  191,
    18921 to 19016 =>  192,
    19017 to 19113 =>  193,
    19114 to 19209 =>  194,
    19210 to 19305 =>  195,
    19306 to 19402 =>  196,
    19403 to 19498 =>  197,
    19499 to 19594 =>  198,
    19595 to 19690 =>  199,
    19691 to 19787 =>  200,
    19788 to 19883 =>  201,
    19884 to 19979 =>  202,
    19980 to 20075 =>  203,
    20076 to 20171 =>  204,
    20172 to 20267 =>  205,
    20268 to 20363 =>  206,
    20364 to 20459 =>  207,
    20460 to 20555 =>  208,
    20556 to 20650 =>  209,
    20651 to 20746 =>  210,
    20747 to 20842 =>  211,
    20843 to 20938 =>  212,
    20939 to 21033 =>  213,
    21034 to 21129 =>  214,
    21130 to 21224 =>  215,
    21225 to 21320 =>  216,
    21321 to 21415 =>  217,
    21416 to 21511 =>  218,
    21512 to 21606 =>  219,
    21607 to 21702 =>  220,
    21703 to 21797 =>  221,
    21798 to 21892 =>  222,
    21893 to 21988 =>  223,
    21989 to 22083 =>  224,
    22084 to 22178 =>  225,
    22179 to 22273 =>  226,
    22274 to 22368 =>  227,
    22369 to 22463 =>  228,
    22464 to 22558 =>  229,
    22559 to 22653 =>  230,
    22654 to 22748 =>  231,
    22749 to 22843 =>  232,
    22844 to 22938 =>  233,
    22939 to 23033 =>  234,
    23034 to 23128 =>  235,
    23129 to 23222 =>  236,
    23223 to 23317 =>  237,
    23318 to 23412 =>  238,
    23413 to 23506 =>  239,
    23507 to 23601 =>  240,
    23602 to 23695 =>  241,
    23696 to 23790 =>  242,
    23791 to 23884 =>  243,
    23885 to 23979 =>  244,
    23980 to 24073 =>  245,
    24074 to 24167 =>  246,
    24168 to 24261 =>  247,
    24262 to 24356 =>  248,
    24357 to 24450 =>  249,
    24451 to 24544 =>  250,
    24545 to 24638 =>  251,
    24639 to 24732 =>  252,
    24733 to 24826 =>  253,
    24827 to 24920 =>  254,
    24921 to 25014 =>  255,
    25015 to 25108 =>  256,
    25109 to 25201 =>  257,
    25202 to 25295 =>  258,
    25296 to 25389 =>  259,
    25390 to 25483 =>  260,
    25484 to 25576 =>  261,
    25577 to 25670 =>  262,
    25671 to 25763 =>  263,
    25764 to 25857 =>  264,
    25858 to 25950 =>  265,
    25951 to 26044 =>  266,
    26045 to 26137 =>  267,
    26138 to 26230 =>  268,
    26231 to 26324 =>  269,
    26325 to 26417 =>  270,
    26418 to 26510 =>  271,
    26511 to 26603 =>  272,
    26604 to 26696 =>  273,
    26697 to 26789 =>  274,
    26790 to 26882 =>  275,
    26883 to 26975 =>  276,
    26976 to 27068 =>  277,
    27069 to 27161 =>  278,
    27162 to 27253 =>  279,
    27254 to 27346 =>  280,
    27347 to 27439 =>  281,
    27440 to 27532 =>  282,
    27533 to 27624 =>  283,
    27625 to 27717 =>  284,
    27718 to 27809 =>  285,
    27810 to 27902 =>  286,
    27903 to 27994 =>  287,
    27995 to 28086 =>  288,
    28087 to 28179 =>  289,
    28180 to 28271 =>  290,
    28272 to 28363 =>  291,
    28364 to 28455 =>  292,
    28456 to 28547 =>  293,
    28548 to 28639 =>  294,
    28640 to 28731 =>  295,
    28732 to 28823 =>  296,
    28824 to 28915 =>  297,
    28916 to 29007 =>  298,
    29008 to 29099 =>  299,
    29100 to 29191 =>  300,
    29192 to 29282 =>  301,
    29283 to 29374 =>  302,
    29375 to 29465 =>  303,
    29466 to 29557 =>  304,
    29558 to 29648 =>  305,
    29649 to 29740 =>  306,
    29741 to 29831 =>  307,
    29832 to 29923 =>  308,
    29924 to 30014 =>  309,
    30015 to 30105 =>  310,
    30106 to 30196 =>  311,
    30197 to 30287 =>  312,
    30288 to 30379 =>  313,
    30380 to 30470 =>  314,
    30471 to 30561 =>  315,
    30562 to 30651 =>  316,
    30652 to 30742 =>  317,
    30743 to 30833 =>  318,
    30834 to 30924 =>  319,
    30925 to 31015 =>  320,
    31016 to 31105 =>  321,
    31106 to 31196 =>  322,
    31197 to 31286 =>  323,
    31287 to 31377 =>  324,
    31378 to 31467 =>  325,
    31468 to 31558 =>  326,
    31559 to 31648 =>  327,
    31649 to 31738 =>  328,
    31739 to 31829 =>  329,
    31830 to 31919 =>  330,
    31920 to 32009 =>  331,
    32010 to 32099 =>  332,
    32100 to 32189 =>  333,
    32190 to 32279 =>  334,
    32280 to 32369 =>  335,
    32370 to 32459 =>  336,
    32460 to 32549 =>  337,
    32550 to 32638 =>  338,
    32639 to 32728 =>  339,
    32729 to 32818 =>  340,
    32819 to 32907 =>  341,
    32908 to 32997 =>  342,
    32998 to 33086 =>  343,
    33087 to 33176 =>  344,
    33177 to 33265 =>  345,
    33266 to 33354 =>  346,
    33355 to 33444 =>  347,
    33445 to 33533 =>  348,
    33534 to 33622 =>  349,
    33623 to 33711 =>  350,
    33712 to 33800 =>  351,
    33801 to 33889 =>  352,
    33890 to 33978 =>  353,
    33979 to 34067 =>  354,
    34068 to 34156 =>  355,
    34157 to 34244 =>  356,
    34245 to 34333 =>  357,
    34334 to 34422 =>  358,
    34423 to 34510 =>  359,
    34511 to 34599 =>  360,
    34600 to 34687 =>  361,
    34688 to 34776 =>  362,
    34777 to 34864 =>  363,
    34865 to 34952 =>  364,
    34953 to 35041 =>  365,
    35042 to 35129 =>  366,
    35130 to 35217 =>  367,
    35218 to 35305 =>  368,
    35306 to 35393 =>  369,
    35394 to 35481 =>  370,
    35482 to 35569 =>  371,
    35570 to 35657 =>  372,
    35658 to 35744 =>  373,
    35745 to 35832 =>  374,
    35833 to 35920 =>  375,
    35921 to 36008 =>  376,
    36009 to 36095 =>  377,
    36096 to 36183 =>  378,
    36184 to 36270 =>  379,
    36271 to 36357 =>  380,
    36358 to 36445 =>  381,
    36446 to 36532 =>  382,
    36533 to 36619 =>  383,
    36620 to 36706 =>  384,
    36707 to 36793 =>  385,
    36794 to 36880 =>  386,
    36881 to 36967 =>  387,
    36968 to 37054 =>  388,
    37055 to 37141 =>  389,
    37142 to 37228 =>  390,
    37229 to 37315 =>  391,
    37316 to 37401 =>  392,
    37402 to 37488 =>  393,
    37489 to 37575 =>  394,
    37576 to 37661 =>  395,
    37662 to 37748 =>  396,
    37749 to 37834 =>  397,
    37835 to 37920 =>  398,
    37921 to 38007 =>  399,
    38008 to 38093 =>  400,
    38094 to 38179 =>  401,
    38180 to 38265 =>  402,
    38266 to 38351 =>  403,
    38352 to 38437 =>  404,
    38438 to 38523 =>  405,
    38524 to 38609 =>  406,
    38610 to 38695 =>  407,
    38696 to 38780 =>  408,
    38781 to 38866 =>  409,
    38867 to 38952 =>  410,
    38953 to 39037 =>  411,
    39038 to 39123 =>  412,
    39124 to 39208 =>  413,
    39209 to 39293 =>  414,
    39294 to 39379 =>  415,
    39380 to 39464 =>  416,
    39465 to 39549 =>  417,
    39550 to 39634 =>  418,
    39635 to 39719 =>  419,
    39720 to 39804 =>  420,
    39805 to 39889 =>  421,
    39890 to 39974 =>  422,
    39975 to 40059 =>  423,
    40060 to 40144 =>  424,
    40145 to 40228 =>  425,
    40229 to 40313 =>  426,
    40314 to 40398 =>  427,
    40399 to 40482 =>  428,
    40483 to 40567 =>  429,
    40568 to 40651 =>  430,
    40652 to 40735 =>  431,
    40736 to 40820 =>  432,
    40821 to 40904 =>  433,
    40905 to 40988 =>  434,
    40989 to 41072 =>  435,
    41073 to 41156 =>  436,
    41157 to 41240 =>  437,
    41241 to 41324 =>  438,
    41325 to 41408 =>  439,
    41409 to 41492 =>  440,
    41493 to 41575 =>  441,
    41576 to 41659 =>  442,
    41660 to 41743 =>  443,
    41744 to 41826 =>  444,
    41827 to 41910 =>  445,
    41911 to 41993 =>  446,
    41994 to 42076 =>  447,
    42077 to 42160 =>  448,
    42161 to 42243 =>  449,
    42244 to 42326 =>  450,
    42327 to 42409 =>  451,
    42410 to 42492 =>  452,
    42493 to 42575 =>  453,
    42576 to 42658 =>  454,
    42659 to 42741 =>  455,
    42742 to 42824 =>  456,
    42825 to 42906 =>  457,
    42907 to 42989 =>  458,
    42990 to 43072 =>  459,
    43073 to 43154 =>  460,
    43155 to 43237 =>  461,
    43238 to 43319 =>  462,
    43320 to 43401 =>  463,
    43402 to 43484 =>  464,
    43485 to 43566 =>  465,
    43567 to 43648 =>  466,
    43649 to 43730 =>  467,
    43731 to 43812 =>  468,
    43813 to 43894 =>  469,
    43895 to 43976 =>  470,
    43977 to 44058 =>  471,
    44059 to 44140 =>  472,
    44141 to 44221 =>  473,
    44222 to 44303 =>  474,
    44304 to 44385 =>  475,
    44386 to 44466 =>  476,
    44467 to 44548 =>  477,
    44549 to 44629 =>  478,
    44630 to 44710 =>  479,
    44711 to 44792 =>  480,
    44793 to 44873 =>  481,
    44874 to 44954 =>  482,
    44955 to 45035 =>  483,
    45036 to 45116 =>  484,
    45117 to 45197 =>  485,
    45198 to 45278 =>  486,
    45279 to 45359 =>  487,
    45360 to 45440 =>  488,
    45441 to 45520 =>  489,
    45521 to 45601 =>  490,
    45602 to 45681 =>  491,
    45682 to 45762 =>  492,
    45763 to 45842 =>  493,
    45843 to 45923 =>  494,
    45924 to 46003 =>  495,
    46004 to 46083 =>  496,
    46084 to 46164 =>  497,
    46165 to 46244 =>  498,
    46245 to 46324 =>  499,
    46325 to 46404 =>  500,
    46405 to 46484 =>  501,
    46485 to 46564 =>  502,
    46565 to 46643 =>  503,
    46644 to 46723 =>  504,
    46724 to 46803 =>  505,
    46804 to 46882 =>  506,
    46883 to 46962 =>  507,
    46963 to 47041 =>  508,
    47042 to 47121 =>  509,
    47122 to 47200 =>  510,
    47201 to 47280 =>  511,
    47281 to 47359 =>  512,
    47360 to 47438 =>  513,
    47439 to 47517 =>  514,
    47518 to 47596 =>  515,
    47597 to 47675 =>  516,
    47676 to 47754 =>  517,
    47755 to 47833 =>  518,
    47834 to 47912 =>  519,
    47913 to 47990 =>  520,
    47991 to 48069 =>  521,
    48070 to 48148 =>  522,
    48149 to 48226 =>  523,
    48227 to 48304 =>  524,
    48305 to 48383 =>  525,
    48384 to 48461 =>  526,
    48462 to 48539 =>  527,
    48540 to 48618 =>  528,
    48619 to 48696 =>  529,
    48697 to 48774 =>  530,
    48775 to 48852 =>  531,
    48853 to 48930 =>  532,
    48931 to 49008 =>  533,
    49009 to 49086 =>  534,
    49087 to 49163 =>  535,
    49164 to 49241 =>  536,
    49242 to 49319 =>  537,
    49320 to 49396 =>  538,
    49397 to 49474 =>  539,
    49475 to 49551 =>  540,
    49552 to 49628 =>  541,
    49629 to 49706 =>  542,
    49707 to 49783 =>  543,
    49784 to 49860 =>  544,
    49861 to 49937 =>  545,
    49938 to 50014 =>  546,
    50015 to 50091 =>  547,
    50092 to 50168 =>  548,
    50169 to 50245 =>  549,
    50246 to 50322 =>  550,
    50323 to 50398 =>  551,
    50399 to 50475 =>  552,
    50476 to 50552 =>  553,
    50553 to 50628 =>  554,
    50629 to 50705 =>  555,
    50706 to 50781 =>  556,
    50782 to 50857 =>  557,
    50858 to 50934 =>  558,
    50935 to 51010 =>  559,
    51011 to 51086 =>  560,
    51087 to 51162 =>  561,
    51163 to 51238 =>  562,
    51239 to 51314 =>  563,
    51315 to 51390 =>  564,
    51391 to 51466 =>  565,
    51467 to 51541 =>  566,
    51542 to 51617 =>  567,
    51618 to 51693 =>  568,
    51694 to 51768 =>  569,
    51769 to 51844 =>  570,
    51845 to 51919 =>  571,
    51920 to 51994 =>  572,
    51995 to 52070 =>  573,
    52071 to 52145 =>  574,
    52146 to 52220 =>  575,
    52221 to 52295 =>  576,
    52296 to 52370 =>  577,
    52371 to 52445 =>  578,
    52446 to 52520 =>  579,
    52521 to 52595 =>  580,
    52596 to 52670 =>  581,
    52671 to 52744 =>  582,
    52745 to 52819 =>  583,
    52820 to 52893 =>  584,
    52894 to 52968 =>  585,
    52969 to 53042 =>  586,
    53043 to 53117 =>  587,
    53118 to 53191 =>  588,
    53192 to 53265 =>  589,
    53266 to 53339 =>  590,
    53340 to 53414 =>  591,
    53415 to 53488 =>  592,
    53489 to 53562 =>  593,
    53563 to 53636 =>  594,
    53637 to 53709 =>  595,
    53710 to 53783 =>  596,
    53784 to 53857 =>  597,
    53858 to 53931 =>  598,
    53932 to 54004 =>  599,
    54005 to 54078 =>  600,
    54079 to 54151 =>  601,
    54152 to 54225 =>  602,
    54226 to 54298 =>  603,
    54299 to 54371 =>  604,
    54372 to 54444 =>  605,
    54445 to 54518 =>  606,
    54519 to 54591 =>  607,
    54592 to 54664 =>  608,
    54665 to 54737 =>  609,
    54738 to 54809 =>  610,
    54810 to 54882 =>  611,
    54883 to 54955 =>  612,
    54956 to 55028 =>  613,
    55029 to 55100 =>  614,
    55101 to 55173 =>  615,
    55174 to 55245 =>  616,
    55246 to 55318 =>  617,
    55319 to 55390 =>  618,
    55391 to 55462 =>  619,
    55463 to 55535 =>  620,
    55536 to 55607 =>  621,
    55608 to 55679 =>  622,
    55680 to 55751 =>  623,
    55752 to 55823 =>  624,
    55824 to 55895 =>  625,
    55896 to 55967 =>  626,
    55968 to 56038 =>  627,
    56039 to 56110 =>  628,
    56111 to 56182 =>  629,
    56183 to 56253 =>  630,
    56254 to 56325 =>  631,
    56326 to 56396 =>  632,
    56397 to 56468 =>  633,
    56469 to 56539 =>  634,
    56540 to 56610 =>  635,
    56611 to 56682 =>  636,
    56683 to 56753 =>  637,
    56754 to 56824 =>  638,
    56825 to 56895 =>  639,
    56896 to 56966 =>  640,
    56967 to 57037 =>  641,
    57038 to 57107 =>  642,
    57108 to 57178 =>  643,
    57179 to 57249 =>  644,
    57250 to 57320 =>  645,
    57321 to 57390 =>  646,
    57391 to 57461 =>  647,
    57462 to 57531 =>  648,
    57532 to 57601 =>  649,
    57602 to 57672 =>  650,
    57673 to 57742 =>  651,
    57743 to 57812 =>  652,
    57813 to 57882 =>  653,
    57883 to 57952 =>  654,
    57953 to 58022 =>  655,
    58023 to 58092 =>  656,
    58093 to 58162 =>  657,
    58163 to 58232 =>  658,
    58233 to 58301 =>  659,
    58302 to 58371 =>  660,
    58372 to 58441 =>  661,
    58442 to 58510 =>  662,
    58511 to 58580 =>  663,
    58581 to 58649 =>  664,
    58650 to 58718 =>  665,
    58719 to 58788 =>  666,
    58789 to 58857 =>  667,
    58858 to 58926 =>  668,
    58927 to 58995 =>  669,
    58996 to 59064 =>  670,
    59065 to 59133 =>  671,
    59134 to 59202 =>  672,
    59203 to 59271 =>  673,
    59272 to 59340 =>  674,
    59341 to 59408 =>  675,
    59409 to 59477 =>  676,
    59478 to 59546 =>  677,
    59547 to 59614 =>  678,
    59615 to 59682 =>  679,
    59683 to 59751 =>  680,
    59752 to 59819 =>  681,
    59820 to 59887 =>  682,
    59888 to 59956 =>  683,
    59957 to 60024 =>  684,
    60025 to 60092 =>  685,
    60093 to 60160 =>  686,
    60161 to 60228 =>  687,
    60229 to 60296 =>  688,
    60297 to 60363 =>  689,
    60364 to 60431 =>  690,
    60432 to 60499 =>  691,
    60500 to 60566 =>  692,
    60567 to 60634 =>  693,
    60635 to 60702 =>  694,
    60703 to 60769 =>  695,
    60770 to 60836 =>  696,
    60837 to 60904 =>  697,
    60905 to 60971 =>  698,
    60972 to 61038 =>  699,
    61039 to 61105 =>  700,
    61106 to 61172 =>  701,
    61173 to 61239 =>  702,
    61240 to 61306 =>  703,
    61307 to 61373 =>  704,
    61374 to 61440 =>  705,
    61441 to 61506 =>  706,
    61507 to 61573 =>  707,
    61574 to 61640 =>  708,
    61641 to 61706 =>  709,
    61707 to 61773 =>  710,
    61774 to 61839 =>  711,
    61840 to 61906 =>  712,
    61907 to 61972 =>  713,
    61973 to 62038 =>  714,
    62039 to 62104 =>  715,
    62105 to 62170 =>  716,
    62171 to 62236 =>  717,
    62237 to 62302 =>  718,
    62303 to 62368 =>  719,
    62369 to 62434 =>  720,
    62435 to 62500 =>  721,
    62501 to 62566 =>  722,
    62567 to 62631 =>  723,
    62632 to 62697 =>  724,
    62698 to 62763 =>  725,
    62764 to 62828 =>  726,
    62829 to 62893 =>  727,
    62894 to 62959 =>  728,
    62960 to 63024 =>  729,
    63025 to 63089 =>  730,
    63090 to 63155 =>  731,
    63156 to 63220 =>  732,
    63221 to 63285 =>  733,
    63286 to 63350 =>  734,
    63351 to 63415 =>  735,
    63416 to 63479 =>  736,
    63480 to 63544 =>  737,
    63545 to 63609 =>  738,
    63610 to 63674 =>  739,
    63675 to 63738 =>  740,
    63739 to 63803 =>  741,
    63804 to 63867 =>  742,
    63868 to 63932 =>  743,
    63933 to 63996 =>  744,
    63997 to 64060 =>  745,
    64061 to 64125 =>  746,
    64126 to 64189 =>  747,
    64190 to 64253 =>  748,
    64254 to 64317 =>  749,
    64318 to 64381 =>  750,
    64382 to 64445 =>  751,
    64446 to 64509 =>  752,
    64510 to 64573 =>  753,
    64574 to 64636 =>  754,
    64637 to 64700 =>  755,
    64701 to 64764 =>  756,
    64765 to 64827 =>  757,
    64828 to 64891 =>  758,
    64892 to 64954 =>  759,
    64955 to 65018 =>  760,
    65019 to 65081 =>  761,
    65082 to 65144 =>  762,
    65145 to 65208 =>  763,
    65209 to 65271 =>  764,
    65272 to 65334 =>  765,
    65335 to 65397 =>  766,
    65398 to 65460 =>  767,
    65461 to 65523 =>  768,
    65524 to 65585 =>  769,
    65586 to 65648 =>  770,
    65649 to 65711 =>  771,
    65712 to 65774 =>  772,
    65775 to 65836 =>  773,
    65837 to 65899 =>  774,
    65900 to 65961 =>  775,
    65962 to 66024 =>  776,
    66025 to 66086 =>  777,
    66087 to 66148 =>  778,
    66149 to 66211 =>  779,
    66212 to 66273 =>  780,
    66274 to 66335 =>  781,
    66336 to 66397 =>  782,
    66398 to 66459 =>  783,
    66460 to 66521 =>  784,
    66522 to 66583 =>  785,
    66584 to 66644 =>  786,
    66645 to 66706 =>  787,
    66707 to 66768 =>  788,
    66769 to 66830 =>  789,
    66831 to 66891 =>  790,
    66892 to 66953 =>  791,
    66954 to 67014 =>  792,
    67015 to 67075 =>  793,
    67076 to 67137 =>  794,
    67138 to 67198 =>  795,
    67199 to 67259 =>  796,
    67260 to 67320 =>  797,
    67321 to 67382 =>  798,
    67383 to 67443 =>  799,
    67444 to 67504 =>  800,
    67505 to 67564 =>  801,
    67565 to 67625 =>  802,
    67626 to 67686 =>  803,
    67687 to 67747 =>  804,
    67748 to 67808 =>  805,
    67809 to 67868 =>  806,
    67869 to 67929 =>  807,
    67930 to 67989 =>  808,
    67990 to 68050 =>  809,
    68051 to 68110 =>  810,
    68111 to 68170 =>  811,
    68171 to 68231 =>  812,
    68232 to 68291 =>  813,
    68292 to 68351 =>  814,
    68352 to 68411 =>  815,
    68412 to 68471 =>  816,
    68472 to 68531 =>  817,
    68532 to 68591 =>  818,
    68592 to 68651 =>  819,
    68652 to 68711 =>  820,
    68712 to 68770 =>  821,
    68771 to 68830 =>  822,
    68831 to 68890 =>  823,
    68891 to 68949 =>  824,
    68950 to 69009 =>  825,
    69010 to 69068 =>  826,
    69069 to 69128 =>  827,
    69129 to 69187 =>  828,
    69188 to 69246 =>  829,
    69247 to 69305 =>  830,
    69306 to 69365 =>  831,
    69366 to 69424 =>  832,
    69425 to 69483 =>  833,
    69484 to 69542 =>  834,
    69543 to 69601 =>  835,
    69602 to 69659 =>  836,
    69660 to 69718 =>  837,
    69719 to 69777 =>  838,
    69778 to 69836 =>  839,
    69837 to 69894 =>  840,
    69895 to 69953 =>  841,
    69954 to 70011 =>  842,
    70012 to 70070 =>  843,
    70071 to 70128 =>  844,
    70129 to 70187 =>  845,
    70188 to 70245 =>  846,
    70246 to 70303 =>  847,
    70304 to 70361 =>  848,
    70362 to 70419 =>  849,
    70420 to 70477 =>  850,
    70478 to 70535 =>  851,
    70536 to 70593 =>  852,
    70594 to 70651 =>  853,
    70652 to 70709 =>  854,
    70710 to 70767 =>  855,
    70768 to 70825 =>  856,
    70826 to 70882 =>  857,
    70883 to 70940 =>  858,
    70941 to 70997 =>  859,
    70998 to 71055 =>  860,
    71056 to 71112 =>  861,
    71113 to 71170 =>  862,
    71171 to 71227 =>  863,
    71228 to 71284 =>  864,
    71285 to 71341 =>  865,
    71342 to 71399 =>  866,
    71400 to 71456 =>  867,
    71457 to 71513 =>  868,
    71514 to 71570 =>  869,
    71571 to 71627 =>  870,
    71628 to 71683 =>  871,
    71684 to 71740 =>  872,
    71741 to 71797 =>  873,
    71798 to 71854 =>  874,
    71855 to 71910 =>  875,
    71911 to 71967 =>  876,
    71968 to 72023 =>  877,
    72024 to 72080 =>  878,
    72081 to 72136 =>  879,
    72137 to 72193 =>  880,
    72194 to 72249 =>  881,
    72250 to 72305 =>  882,
    72306 to 72361 =>  883,
    72362 to 72418 =>  884,
    72419 to 72474 =>  885,
    72475 to 72530 =>  886,
    72531 to 72586 =>  887,
    72587 to 72641 =>  888,
    72642 to 72697 =>  889,
    72698 to 72753 =>  890,
    72754 to 72809 =>  891,
    72810 to 72865 =>  892,
    72866 to 72920 =>  893,
    72921 to 72976 =>  894,
    72977 to 73031 =>  895,
    73032 to 73087 =>  896,
    73088 to 73142 =>  897,
    73143 to 73198 =>  898,
    73199 to 73253 =>  899,
    73254 to 73308 =>  900,
    73309 to 73363 =>  901,
    73364 to 73418 =>  902,
    73419 to 73474 =>  903,
    73475 to 73529 =>  904,
    73530 to 73584 =>  905,
    73585 to 73638 =>  906,
    73639 to 73693 =>  907,
    73694 to 73748 =>  908,
    73749 to 73803 =>  909,
    73804 to 73858 =>  910,
    73859 to 73912 =>  911,
    73913 to 73967 =>  912,
    73968 to 74021 =>  913,
    74022 to 74076 =>  914,
    74077 to 74130 =>  915,
    74131 to 74185 =>  916,
    74186 to 74239 =>  917,
    74240 to 74293 =>  918,
    74294 to 74347 =>  919,
    74348 to 74402 =>  920,
    74403 to 74456 =>  921,
    74457 to 74510 =>  922,
    74511 to 74564 =>  923,
    74565 to 74618 =>  924,
    74619 to 74672 =>  925,
    74673 to 74725 =>  926,
    74726 to 74779 =>  927,
    74780 to 74833 =>  928,
    74834 to 74887 =>  929,
    74888 to 74940 =>  930,
    74941 to 74994 =>  931,
    74995 to 75047 =>  932,
    75048 to 75101 =>  933,
    75102 to 75154 =>  934,
    75155 to 75208 =>  935,
    75209 to 75261 =>  936,
    75262 to 75314 =>  937,
    75315 to 75367 =>  938,
    75368 to 75420 =>  939,
    75421 to 75474 =>  940,
    75475 to 75527 =>  941,
    75528 to 75580 =>  942,
    75581 to 75633 =>  943,
    75634 to 75685 =>  944,
    75686 to 75738 =>  945,
    75739 to 75791 =>  946,
    75792 to 75844 =>  947,
    75845 to 75896 =>  948,
    75897 to 75949 =>  949,
    75950 to 76002 =>  950,
    76003 to 76054 =>  951,
    76055 to 76107 =>  952,
    76108 to 76159 =>  953,
    76160 to 76211 =>  954,
    76212 to 76264 =>  955,
    76265 to 76316 =>  956,
    76317 to 76368 =>  957,
    76369 to 76420 =>  958,
    76421 to 76472 =>  959,
    76473 to 76524 =>  960,
    76525 to 76576 =>  961,
    76577 to 76628 =>  962,
    76629 to 76680 =>  963,
    76681 to 76732 =>  964,
    76733 to 76784 =>  965,
    76785 to 76835 =>  966,
    76836 to 76887 =>  967,
    76888 to 76939 =>  968,
    76940 to 76990 =>  969,
    76991 to 77042 =>  970,
    77043 to 77093 =>  971,
    77094 to 77145 =>  972,
    77146 to 77196 =>  973,
    77197 to 77247 =>  974,
    77248 to 77299 =>  975,
    77300 to 77350 =>  976,
    77351 to 77401 =>  977,
    77402 to 77452 =>  978,
    77453 to 77503 =>  979,
    77504 to 77554 =>  980,
    77555 to 77605 =>  981,
    77606 to 77656 =>  982,
    77657 to 77707 =>  983,
    77708 to 77758 =>  984,
    77759 to 77809 =>  985,
    77810 to 77859 =>  986,
    77860 to 77910 =>  987,
    77911 to 77960 =>  988,
    77961 to 78011 =>  989,
    78012 to 78062 =>  990,
    78063 to 78112 =>  991,
    78113 to 78162 =>  992,
    78163 to 78213 =>  993,
    78214 to 78263 =>  994,
    78264 to 78313 =>  995,
    78314 to 78364 =>  996,
    78365 to 78414 =>  997,
    78415 to 78464 =>  998,
    78465 to 78514 =>  999,
    78515 to 78564 => 1000,
    78565 to 78614 => 1001,
    78615 to 78664 => 1002,
    78665 to 78714 => 1003,
    78715 to 78763 => 1004,
    78764 to 78813 => 1005,
    78814 to 78863 => 1006,
    78864 to 78912 => 1007,
    78913 to 78962 => 1008,
    78963 to 79012 => 1009,
    79013 to 79061 => 1010,
    79062 to 79111 => 1011,
    79112 to 79160 => 1012,
    79161 to 79209 => 1013,
    79210 to 79259 => 1014,
    79260 to 79308 => 1015,
    79309 to 79357 => 1016,
    79358 to 79406 => 1017,
    79407 to 79455 => 1018,
    79456 to 79504 => 1019,
    79505 to 79553 => 1020,
    79554 to 79602 => 1021,
    79603 to 79651 => 1022,
    79652 to 79700 => 1023,
    79701 to 79749 => 1024,
    79750 to 79798 => 1025,
    79799 to 79846 => 1026,
    79847 to 79895 => 1027,
    79896 to 79944 => 1028,
    79945 to 79992 => 1029,
    79993 to 80041 => 1030,
    80042 to 80089 => 1031,
    80090 to 80138 => 1032,
    80139 to 80186 => 1033,
    80187 to 80234 => 1034,
    80235 to 80283 => 1035,
    80284 to 80331 => 1036,
    80332 to 80379 => 1037,
    80380 to 80427 => 1038,
    80428 to 80475 => 1039,
    80476 to 80523 => 1040,
    80524 to 80571 => 1041,
    80572 to 80619 => 1042,
    80620 to 80667 => 1043,
    80668 to 80715 => 1044,
    80716 to 80763 => 1045,
    80764 to 80811 => 1046,
    80812 to 80858 => 1047,
    80859 to 80906 => 1048,
    80907 to 80954 => 1049,
    80955 to 81001 => 1050,
    81002 to 81049 => 1051,
    81050 to 81096 => 1052,
    81097 to 81144 => 1053,
    81145 to 81191 => 1054,
    81192 to 81238 => 1055,
    81239 to 81286 => 1056,
    81287 to 81333 => 1057,
    81334 to 81380 => 1058,
    81381 to 81427 => 1059,
    81428 to 81474 => 1060,
    81475 to 81521 => 1061,
    81522 to 81568 => 1062,
    81569 to 81615 => 1063,
    81616 to 81662 => 1064,
    81663 to 81709 => 1065,
    81710 to 81756 => 1066,
    81757 to 81802 => 1067,
    81803 to 81849 => 1068,
    81850 to 81896 => 1069,
    81897 to 81942 => 1070,
    81943 to 81989 => 1071,
    81990 to 82036 => 1072,
    82037 to 82082 => 1073,
    82083 to 82128 => 1074,
    82129 to 82175 => 1075,
    82176 to 82221 => 1076,
    82222 to 82268 => 1077,
    82269 to 82314 => 1078,
    82315 to 82360 => 1079,
    82361 to 82406 => 1080,
    82407 to 82452 => 1081,
    82453 to 82498 => 1082,
    82499 to 82544 => 1083,
    82545 to 82590 => 1084,
    82591 to 82636 => 1085,
    82637 to 82682 => 1086,
    82683 to 82728 => 1087,
    82729 to 82774 => 1088,
    82775 to 82820 => 1089,
    82821 to 82865 => 1090,
    82866 to 82911 => 1091,
    82912 to 82956 => 1092,
    82957 to 83002 => 1093,
    83003 to 83048 => 1094,
    83049 to 83093 => 1095,
    83094 to 83138 => 1096,
    83139 to 83184 => 1097,
    83185 to 83229 => 1098,
    83230 to 83274 => 1099,
    83275 to 83320 => 1100,
    83321 to 83365 => 1101,
    83366 to 83410 => 1102,
    83411 to 83455 => 1103,
    83456 to 83500 => 1104,
    83501 to 83545 => 1105,
    83546 to 83590 => 1106,
    83591 to 83635 => 1107,
    83636 to 83680 => 1108,
    83681 to 83725 => 1109,
    83726 to 83770 => 1110,
    83771 to 83815 => 1111,
    83816 to 83859 => 1112,
    83860 to 83904 => 1113,
    83905 to 83949 => 1114,
    83950 to 83993 => 1115,
    83994 to 84038 => 1116,
    84039 to 84082 => 1117,
    84083 to 84127 => 1118,
    84128 to 84171 => 1119,
    84172 to 84215 => 1120,
    84216 to 84260 => 1121,
    84261 to 84304 => 1122,
    84305 to 84348 => 1123,
    84349 to 84392 => 1124,
    84393 to 84436 => 1125,
    84437 to 84481 => 1126,
    84482 to 84525 => 1127,
    84526 to 84569 => 1128,
    84570 to 84613 => 1129,
    84614 to 84656 => 1130,
    84657 to 84700 => 1131,
    84701 to 84744 => 1132,
    84745 to 84788 => 1133,
    84789 to 84832 => 1134,
    84833 to 84875 => 1135,
    84876 to 84919 => 1136,
    84920 to 84963 => 1137,
    84964 to 85006 => 1138,
    85007 to 85050 => 1139,
    85051 to 85093 => 1140,
    85094 to 85137 => 1141,
    85138 to 85180 => 1142,
    85181 to 85223 => 1143,
    85224 to 85267 => 1144,
    85268 to 85310 => 1145,
    85311 to 85353 => 1146,
    85354 to 85396 => 1147,
    85397 to 85440 => 1148,
    85441 to 85483 => 1149,
    85484 to 85526 => 1150,
    85527 to 85569 => 1151,
    85570 to 85612 => 1152,
    85613 to 85655 => 1153,
    85656 to 85698 => 1154,
    85699 to 85740 => 1155,
    85741 to 85783 => 1156,
    85784 to 85826 => 1157,
    85827 to 85869 => 1158,
    85870 to 85911 => 1159,
    85912 to 85954 => 1160,
    85955 to 85997 => 1161,
    85998 to 86039 => 1162,
    86040 to 86082 => 1163,
    86083 to 86124 => 1164,
    86125 to 86167 => 1165,
    86168 to 86209 => 1166,
    86210 to 86251 => 1167,
    86252 to 86294 => 1168,
    86295 to 86336 => 1169,
    86337 to 86378 => 1170,
    86379 to 86420 => 1171,
    86421 to 86462 => 1172,
    86463 to 86504 => 1173,
    86505 to 86546 => 1174,
    86547 to 86588 => 1175,
    86589 to 86630 => 1176,
    86631 to 86672 => 1177,
    86673 to 86714 => 1178,
    86715 to 86756 => 1179,
    86757 to 86798 => 1180,
    86799 to 86840 => 1181,
    86841 to 86881 => 1182,
    86882 to 86923 => 1183,
    86924 to 86965 => 1184,
    86966 to 87006 => 1185,
    87007 to 87048 => 1186,
    87049 to 87089 => 1187,
    87090 to 87131 => 1188,
    87132 to 87172 => 1189,
    87173 to 87214 => 1190,
    87215 to 87255 => 1191,
    87256 to 87296 => 1192,
    87297 to 87338 => 1193,
    87339 to 87379 => 1194,
    87380 to 87420 => 1195,
    87421 to 87461 => 1196,
    87462 to 87502 => 1197,
    87503 to 87543 => 1198,
    87544 to 87584 => 1199,
    87585 to 87625 => 1200,
    87626 to 87666 => 1201,
    87667 to 87707 => 1202,
    87708 to 87748 => 1203,
    87749 to 87789 => 1204,
    87790 to 87830 => 1205,
    87831 to 87870 => 1206,
    87871 to 87911 => 1207,
    87912 to 87952 => 1208,
    87953 to 87992 => 1209,
    87993 to 88033 => 1210,
    88034 to 88073 => 1211,
    88074 to 88114 => 1212,
    88115 to 88154 => 1213,
    88155 to 88195 => 1214,
    88196 to 88235 => 1215,
    88236 to 88276 => 1216,
    88277 to 88316 => 1217,
    88317 to 88356 => 1218,
    88357 to 88396 => 1219,
    88397 to 88437 => 1220,
    88438 to 88477 => 1221,
    88478 to 88517 => 1222,
    88518 to 88557 => 1223,
    88558 to 88597 => 1224,
    88598 to 88637 => 1225,
    88638 to 88677 => 1226,
    88678 to 88717 => 1227,
    88718 to 88757 => 1228,
    88758 to 88796 => 1229,
    88797 to 88836 => 1230,
    88837 to 88876 => 1231,
    88877 to 88916 => 1232,
    88917 to 88955 => 1233,
    88956 to 88995 => 1234,
    88996 to 89035 => 1235,
    89036 to 89074 => 1236,
    89075 to 89114 => 1237,
    89115 to 89153 => 1238,
    89154 to 89193 => 1239,
    89194 to 89232 => 1240,
    89233 to 89271 => 1241,
    89272 to 89311 => 1242,
    89312 to 89350 => 1243,
    89351 to 89389 => 1244,
    89390 to 89429 => 1245,
    89430 to 89468 => 1246,
    89469 to 89507 => 1247,
    89508 to 89546 => 1248,
    89547 to 89585 => 1249,
    89586 to 89624 => 1250,
    89625 to 89663 => 1251,
    89664 to 89702 => 1252,
    89703 to 89741 => 1253,
    89742 to 89780 => 1254,
    89781 to 89819 => 1255,
    89820 to 89857 => 1256,
    89858 to 89896 => 1257,
    89897 to 89935 => 1258,
    89936 to 89974 => 1259,
    89975 to 90012 => 1260,
    90013 to 90051 => 1261,
    90052 to 90089 => 1262,
    90090 to 90128 => 1263,
    90129 to 90166 => 1264,
    90167 to 90205 => 1265,
    90206 to 90243 => 1266,
    90244 to 90282 => 1267,
    90283 to 90320 => 1268,
    90321 to 90358 => 1269,
    90359 to 90397 => 1270,
    90398 to 90435 => 1271,
    90436 to 90473 => 1272,
    90474 to 90511 => 1273,
    90512 to 90549 => 1274,
    90550 to 90587 => 1275,
    90588 to 90625 => 1276,
    90626 to 90663 => 1277,
    90664 to 90701 => 1278,
    90702 to 90739 => 1279,
    90740 to 90777 => 1280,
    90778 to 90815 => 1281,
    90816 to 90853 => 1282,
    90854 to 90891 => 1283,
    90892 to 90929 => 1284,
    90930 to 90966 => 1285,
    90967 to 91004 => 1286,
    91005 to 91042 => 1287,
    91043 to 91079 => 1288,
    91080 to 91117 => 1289,
    91118 to 91154 => 1290,
    91155 to 91192 => 1291,
    91193 to 91229 => 1292,
    91230 to 91267 => 1293,
    91268 to 91304 => 1294,
    91305 to 91341 => 1295,
    91342 to 91379 => 1296,
    91380 to 91416 => 1297,
    91417 to 91453 => 1298,
    91454 to 91490 => 1299,
    91491 to 91528 => 1300,
    91529 to 91565 => 1301,
    91566 to 91602 => 1302,
    91603 to 91639 => 1303,
    91640 to 91676 => 1304,
    91677 to 91713 => 1305,
    91714 to 91750 => 1306,
    91751 to 91787 => 1307,
    91788 to 91824 => 1308,
    91825 to 91861 => 1309,
    91862 to 91897 => 1310,
    91898 to 91934 => 1311,
    91935 to 91971 => 1312,
    91972 to 92008 => 1313,
    92009 to 92044 => 1314,
    92045 to 92081 => 1315,
    92082 to 92118 => 1316,
    92119 to 92154 => 1317,
    92155 to 92191 => 1318,
    92192 to 92227 => 1319,
    92228 to 92264 => 1320,
    92265 to 92300 => 1321,
    92301 to 92336 => 1322,
    92337 to 92373 => 1323,
    92374 to 92409 => 1324,
    92410 to 92445 => 1325,
    92446 to 92482 => 1326,
    92483 to 92518 => 1327,
    92519 to 92554 => 1328,
    92555 to 92590 => 1329,
    92591 to 92626 => 1330,
    92627 to 92662 => 1331,
    92663 to 92699 => 1332,
    92700 to 92735 => 1333,
    92736 to 92770 => 1334,
    92771 to 92806 => 1335,
    92807 to 92842 => 1336,
    92843 to 92878 => 1337,
    92879 to 92914 => 1338,
    92915 to 92950 => 1339,
    92951 to 92986 => 1340,
    92987 to 93021 => 1341,
    93022 to 93057 => 1342,
    93058 to 93093 => 1343,
    93094 to 93128 => 1344,
    93129 to 93164 => 1345,
    93165 to 93200 => 1346,
    93201 to 93235 => 1347,
    93236 to 93271 => 1348,
    93272 to 93306 => 1349,
    93307 to 93341 => 1350,
    93342 to 93377 => 1351,
    93378 to 93412 => 1352,
    93413 to 93448 => 1353,
    93449 to 93483 => 1354,
    93484 to 93518 => 1355,
    93519 to 93553 => 1356,
    93554 to 93589 => 1357,
    93590 to 93624 => 1358,
    93625 to 93659 => 1359,
    93660 to 93694 => 1360,
    93695 to 93729 => 1361,
    93730 to 93764 => 1362,
    93765 to 93799 => 1363,
    93800 to 93834 => 1364,
    93835 to 93869 => 1365,
    93870 to 93904 => 1366,
    93905 to 93939 => 1367,
    93940 to 93973 => 1368,
    93974 to 94008 => 1369,
    94009 to 94043 => 1370,
    94044 to 94078 => 1371,
    94079 to 94112 => 1372,
    94113 to 94147 => 1373,
    94148 to 94182 => 1374,
    94183 to 94216 => 1375,
    94217 to 94251 => 1376,
    94252 to 94285 => 1377,
    94286 to 94320 => 1378,
    94321 to 94354 => 1379,
    94355 to 94389 => 1380,
    94390 to 94423 => 1381,
    94424 to 94458 => 1382,
    94459 to 94492 => 1383,
    94493 to 94526 => 1384,
    94527 to 94560 => 1385,
    94561 to 94595 => 1386,
    94596 to 94629 => 1387,
    94630 to 94663 => 1388,
    94664 to 94697 => 1389,
    94698 to 94731 => 1390,
    94732 to 94765 => 1391,
    94766 to 94799 => 1392,
    94800 to 94833 => 1393,
    94834 to 94867 => 1394,
    94868 to 94901 => 1395,
    94902 to 94935 => 1396,
    94936 to 94969 => 1397,
    94970 to 95003 => 1398,
    95004 to 95037 => 1399,
    95038 to 95071 => 1400,
    95072 to 95104 => 1401,
    95105 to 95138 => 1402,
    95139 to 95172 => 1403,
    95173 to 95205 => 1404,
    95206 to 95239 => 1405,
    95240 to 95273 => 1406,
    95274 to 95306 => 1407,
    95307 to 95340 => 1408,
    95341 to 95373 => 1409,
    95374 to 95407 => 1410,
    95408 to 95440 => 1411,
    95441 to 95473 => 1412,
    95474 to 95507 => 1413,
    95508 to 95540 => 1414,
    95541 to 95574 => 1415,
    95575 to 95607 => 1416,
    95608 to 95640 => 1417,
    95641 to 95673 => 1418,
    95674 to 95706 => 1419,
    95707 to 95740 => 1420,
    95741 to 95773 => 1421,
    95774 to 95806 => 1422,
    95807 to 95839 => 1423,
    95840 to 95872 => 1424,
    95873 to 95905 => 1425,
    95906 to 95938 => 1426,
    95939 to 95971 => 1427,
    95972 to 96004 => 1428,
    96005 to 96037 => 1429,
    96038 to 96069 => 1430,
    96070 to 96102 => 1431,
    96103 to 96135 => 1432,
    96136 to 96168 => 1433,
    96169 to 96200 => 1434,
    96201 to 96233 => 1435,
    96234 to 96266 => 1436,
    96267 to 96298 => 1437,
    96299 to 96331 => 1438,
    96332 to 96364 => 1439,
    96365 to 96396 => 1440,
    96397 to 96429 => 1441,
    96430 to 96461 => 1442,
    96462 to 96494 => 1443,
    96495 to 96526 => 1444,
    96527 to 96558 => 1445,
    96559 to 96591 => 1446,
    96592 to 96623 => 1447,
    96624 to 96655 => 1448,
    96656 to 96688 => 1449,
    96689 to 96720 => 1450,
    96721 to 96752 => 1451,
    96753 to 96784 => 1452,
    96785 to 96816 => 1453,
    96817 to 96848 => 1454,
    96849 to 96881 => 1455,
    96882 to 96913 => 1456,
    96914 to 96945 => 1457,
    96946 to 96977 => 1458,
    96978 to 97009 => 1459,
    97010 to 97040 => 1460,
    97041 to 97072 => 1461,
    97073 to 97104 => 1462,
    97105 to 97136 => 1463,
    97137 to 97168 => 1464,
    97169 to 97200 => 1465,
    97201 to 97231 => 1466,
    97232 to 97263 => 1467,
    97264 to 97295 => 1468,
    97296 to 97327 => 1469,
    97328 to 97358 => 1470,
    97359 to 97390 => 1471,
    97391 to 97421 => 1472,
    97422 to 97453 => 1473,
    97454 to 97484 => 1474,
    97485 to 97516 => 1475,
    97517 to 97547 => 1476,
    97548 to 97579 => 1477,
    97580 to 97610 => 1478,
    97611 to 97642 => 1479,
    97643 to 97673 => 1480,
    97674 to 97704 => 1481,
    97705 to 97736 => 1482,
    97737 to 97767 => 1483,
    97768 to 97798 => 1484,
    97799 to 97829 => 1485,
    97830 to 97860 => 1486,
    97861 to 97892 => 1487,
    97893 to 97923 => 1488,
    97924 to 97954 => 1489,
    97955 to 97985 => 1490,
    97986 to 98016 => 1491,
    98017 to 98047 => 1492,
    98048 to 98078 => 1493,
    98079 to 98109 => 1494,
    98110 to 98140 => 1495,
    98141 to 98171 => 1496,
    98172 to 98201 => 1497,
    98202 to 98232 => 1498,
    98233 to 98263 => 1499,
    98264 to 98294 => 1500,
    98295 to 98324 => 1501,
    98325 to 98355 => 1502,
    98356 to 98386 => 1503,
    98387 to 98417 => 1504,
    98418 to 98447 => 1505,
    98448 to 98478 => 1506,
    98479 to 98508 => 1507,
    98509 to 98539 => 1508,
    98540 to 98569 => 1509,
    98570 to 98600 => 1510,
    98601 to 98630 => 1511,
    98631 to 98661 => 1512,
    98662 to 98691 => 1513,
    98692 to 98722 => 1514,
    98723 to 98752 => 1515,
    98753 to 98782 => 1516,
    98783 to 98813 => 1517,
    98814 to 98843 => 1518,
    98844 to 98873 => 1519,
    98874 to 98903 => 1520,
    98904 to 98933 => 1521,
    98934 to 98964 => 1522,
    98965 to 98994 => 1523,
    98995 to 99024 => 1524,
    99025 to 99054 => 1525,
    99055 to 99084 => 1526,
    99085 to 99114 => 1527,
    99115 to 99144 => 1528,
    99145 to 99174 => 1529,
    99175 to 99204 => 1530,
    99205 to 99234 => 1531,
    99235 to 99264 => 1532,
    99265 to 99293 => 1533,
    99294 to 99323 => 1534,
    99324 to 99353 => 1535,
    99354 to 99383 => 1536,
    99384 to 99413 => 1537,
    99414 to 99442 => 1538,
    99443 to 99472 => 1539,
    99473 to 99502 => 1540,
    99503 to 99531 => 1541,
    99532 to 99561 => 1542,
    99562 to 99590 => 1543,
    99591 to 99620 => 1544,
    99621 to 99649 => 1545,
    99650 to 99679 => 1546,
    99680 to 99708 => 1547,
    99709 to 99738 => 1548,
    99739 to 99767 => 1549,
    99768 to 99797 => 1550,
    99798 to 99826 => 1551,
    99827 to 99855 => 1552,
    99856 to 99885 => 1553,
    99886 to 99914 => 1554,
    99915 to 99943 => 1555,
    99944 to 99972 => 1556,
    99973 to 100002 => 1557,
    100003 to 100031 => 1558,
    100032 to 100060 => 1559,
    100061 to 100089 => 1560,
    100090 to 100118 => 1561,
    100119 to 100147 => 1562,
    100148 to 100176 => 1563,
    100177 to 100205 => 1564,
    100206 to 100234 => 1565,
    100235 to 100263 => 1566,
    100264 to 100292 => 1567,
    100293 to 100321 => 1568,
    100322 to 100350 => 1569,
    100351 to 100379 => 1570,
    100380 to 100408 => 1571,
    100409 to 100437 => 1572,
    100438 to 100465 => 1573,
    100466 to 100494 => 1574,
    100495 to 100523 => 1575,
    100524 to 100552 => 1576,
    100553 to 100580 => 1577,
    100581 to 100609 => 1578,
    100610 to 100638 => 1579,
    100639 to 100666 => 1580,
    100667 to 100695 => 1581,
    100696 to 100723 => 1582,
    100724 to 100752 => 1583,
    100753 to 100780 => 1584,
    100781 to 100809 => 1585,
    100810 to 100837 => 1586,
    100838 to 100866 => 1587,
    100867 to 100894 => 1588,
    100895 to 100922 => 1589,
    100923 to 100951 => 1590,
    100952 to 100979 => 1591,
    100980 to 101007 => 1592,
    101008 to 101036 => 1593,
    101037 to 101064 => 1594,
    101065 to 101092 => 1595,
    101093 to 101120 => 1596,
    101121 to 101148 => 1597,
    101149 to 101177 => 1598,
    101178 to 101205 => 1599,
    101206 to 101233 => 1600,
    101234 to 101261 => 1601,
    101262 to 101289 => 1602,
    101290 to 101317 => 1603,
    101318 to 101345 => 1604,
    101346 to 101373 => 1605,
    101374 to 101401 => 1606,
    101402 to 101429 => 1607,
    101430 to 101457 => 1608,
    101458 to 101484 => 1609,
    101485 to 101512 => 1610,
    101513 to 101540 => 1611,
    101541 to 101568 => 1612,
    101569 to 101596 => 1613,
    101597 to 101623 => 1614,
    101624 to 101651 => 1615,
    101652 to 101679 => 1616,
    101680 to 101706 => 1617,
    101707 to 101734 => 1618,
    101735 to 101762 => 1619,
    101763 to 101789 => 1620,
    101790 to 101817 => 1621,
    101818 to 101844 => 1622,
    101845 to 101872 => 1623,
    101873 to 101899 => 1624,
    101900 to 101927 => 1625,
    101928 to 101954 => 1626,
    101955 to 101982 => 1627,
    101983 to 102009 => 1628,
    102010 to 102036 => 1629,
    102037 to 102064 => 1630,
    102065 to 102091 => 1631,
    102092 to 102118 => 1632,
    102119 to 102146 => 1633,
    102147 to 102173 => 1634,
    102174 to 102200 => 1635,
    102201 to 102227 => 1636,
    102228 to 102255 => 1637,
    102256 to 102282 => 1638,
    102283 to 102309 => 1639,
    102310 to 102336 => 1640,
    102337 to 102363 => 1641,
    102364 to 102390 => 1642,
    102391 to 102417 => 1643,
    102418 to 102444 => 1644,
    102445 to 102471 => 1645,
    102472 to 102498 => 1646,
    102499 to 102525 => 1647,
    102526 to 102552 => 1648,
    102553 to 102579 => 1649,
    102580 to 102606 => 1650,
    102607 to 102633 => 1651,
    102634 to 102659 => 1652,
    102660 to 102686 => 1653,
    102687 to 102713 => 1654,
    102714 to 102740 => 1655,
    102741 to 102766 => 1656,
    102767 to 102793 => 1657,
    102794 to 102820 => 1658,
    102821 to 102846 => 1659,
    102847 to 102873 => 1660,
    102874 to 102900 => 1661,
    102901 to 102926 => 1662,
    102927 to 102953 => 1663,
    102954 to 102979 => 1664,
    102980 to 103006 => 1665,
    103007 to 103032 => 1666,
    103033 to 103059 => 1667,
    103060 to 103085 => 1668,
    103086 to 103112 => 1669,
    103113 to 103138 => 1670,
    103139 to 103164 => 1671,
    103165 to 103191 => 1672,
    103192 to 103217 => 1673,
    103218 to 103243 => 1674,
    103244 to 103270 => 1675,
    103271 to 103296 => 1676,
    103297 to 103322 => 1677,
    103323 to 103348 => 1678,
    103349 to 103374 => 1679,
    103375 to 103401 => 1680,
    103402 to 103427 => 1681,
    103428 to 103453 => 1682,
    103454 to 103479 => 1683,
    103480 to 103505 => 1684,
    103506 to 103531 => 1685,
    103532 to 103557 => 1686,
    103558 to 103583 => 1687,
    103584 to 103609 => 1688,
    103610 to 103635 => 1689,
    103636 to 103661 => 1690,
    103662 to 103687 => 1691,
    103688 to 103713 => 1692,
    103714 to 103739 => 1693,
    103740 to 103764 => 1694,
    103765 to 103790 => 1695,
    103791 to 103816 => 1696,
    103817 to 103842 => 1697,
    103843 to 103868 => 1698,
    103869 to 103893 => 1699,
    103894 to 103919 => 1700,
    103920 to 103945 => 1701,
    103946 to 103970 => 1702,
    103971 to 103996 => 1703,
    103997 to 104022 => 1704,
    104023 to 104047 => 1705,
    104048 to 104073 => 1706,
    104074 to 104098 => 1707,
    104099 to 104124 => 1708,
    104125 to 104149 => 1709,
    104150 to 104175 => 1710,
    104176 to 104200 => 1711,
    104201 to 104226 => 1712,
    104227 to 104251 => 1713,
    104252 to 104277 => 1714,
    104278 to 104302 => 1715,
    104303 to 104327 => 1716,
    104328 to 104353 => 1717,
    104354 to 104378 => 1718,
    104379 to 104403 => 1719,
    104404 to 104429 => 1720,
    104430 to 104454 => 1721,
    104455 to 104479 => 1722,
    104480 to 104504 => 1723,
    104505 to 104529 => 1724,
    104530 to 104555 => 1725,
    104556 to 104580 => 1726,
    104581 to 104605 => 1727,
    104606 to 104630 => 1728,
    104631 to 104655 => 1729,
    104656 to 104680 => 1730,
    104681 to 104705 => 1731,
    104706 to 104730 => 1732,
    104731 to 104755 => 1733,
    104756 to 104780 => 1734,
    104781 to 104805 => 1735,
    104806 to 104830 => 1736,
    104831 to 104855 => 1737,
    104856 to 104880 => 1738,
    104881 to 104904 => 1739,
    104905 to 104929 => 1740,
    104930 to 104954 => 1741,
    104955 to 104979 => 1742,
    104980 to 105004 => 1743,
    105005 to 105028 => 1744,
    105029 to 105053 => 1745,
    105054 to 105078 => 1746,
    105079 to 105102 => 1747,
    105103 to 105127 => 1748,
    105128 to 105152 => 1749,
    105153 to 105176 => 1750,
    105177 to 105201 => 1751,
    105202 to 105225 => 1752,
    105226 to 105250 => 1753,
    105251 to 105275 => 1754,
    105276 to 105299 => 1755,
    105300 to 105324 => 1756,
    105325 to 105348 => 1757,
    105349 to 105372 => 1758,
    105373 to 105397 => 1759,
    105398 to 105421 => 1760,
    105422 to 105446 => 1761,
    105447 to 105470 => 1762,
    105471 to 105494 => 1763,
    105495 to 105519 => 1764,
    105520 to 105543 => 1765,
    105544 to 105567 => 1766,
    105568 to 105592 => 1767,
    105593 to 105616 => 1768,
    105617 to 105640 => 1769,
    105641 to 105664 => 1770,
    105665 to 105688 => 1771,
    105689 to 105713 => 1772,
    105714 to 105737 => 1773,
    105738 to 105761 => 1774,
    105762 to 105785 => 1775,
    105786 to 105809 => 1776,
    105810 to 105833 => 1777,
    105834 to 105857 => 1778,
    105858 to 105881 => 1779,
    105882 to 105905 => 1780,
    105906 to 105929 => 1781,
    105930 to 105953 => 1782,
    105954 to 105977 => 1783,
    105978 to 106001 => 1784,
    106002 to 106025 => 1785,
    106026 to 106049 => 1786,
    106050 to 106072 => 1787,
    106073 to 106096 => 1788,
    106097 to 106120 => 1789,
    106121 to 106144 => 1790,
    106145 to 106168 => 1791,
    106169 to 106191 => 1792,
    106192 to 106215 => 1793,
    106216 to 106239 => 1794,
    106240 to 106262 => 1795,
    106263 to 106286 => 1796,
    106287 to 106310 => 1797,
    106311 to 106333 => 1798,
    106334 to 106357 => 1799,
    106358 to 106381 => 1800,
    106382 to 106404 => 1801,
    106405 to 106428 => 1802,
    106429 to 106451 => 1803,
    106452 to 106475 => 1804,
    106476 to 106498 => 1805,
    106499 to 106522 => 1806,
    106523 to 106545 => 1807,
    106546 to 106569 => 1808,
    106570 to 106592 => 1809,
    106593 to 106615 => 1810,
    106616 to 106639 => 1811,
    106640 to 106662 => 1812,
    106663 to 106685 => 1813,
    106686 to 106709 => 1814,
    106710 to 106732 => 1815,
    106733 to 106755 => 1816,
    106756 to 106778 => 1817,
    106779 to 106802 => 1818,
    106803 to 106825 => 1819,
    106826 to 106848 => 1820,
    106849 to 106871 => 1821,
    106872 to 106894 => 1822,
    106895 to 106918 => 1823,
    106919 to 106941 => 1824,
    106942 to 106964 => 1825,
    106965 to 106987 => 1826,
    106988 to 107010 => 1827,
    107011 to 107033 => 1828,
    107034 to 107056 => 1829,
    107057 to 107079 => 1830,
    107080 to 107102 => 1831,
    107103 to 107125 => 1832,
    107126 to 107148 => 1833,
    107149 to 107171 => 1834,
    107172 to 107194 => 1835,
    107195 to 107216 => 1836,
    107217 to 107239 => 1837,
    107240 to 107262 => 1838,
    107263 to 107285 => 1839,
    107286 to 107308 => 1840,
    107309 to 107331 => 1841,
    107332 to 107353 => 1842,
    107354 to 107376 => 1843,
    107377 to 107399 => 1844,
    107400 to 107422 => 1845,
    107423 to 107444 => 1846,
    107445 to 107467 => 1847,
    107468 to 107490 => 1848,
    107491 to 107512 => 1849,
    107513 to 107535 => 1850,
    107536 to 107557 => 1851,
    107558 to 107580 => 1852,
    107581 to 107602 => 1853,
    107603 to 107625 => 1854,
    107626 to 107648 => 1855,
    107649 to 107670 => 1856,
    107671 to 107693 => 1857,
    107694 to 107715 => 1858,
    107716 to 107737 => 1859,
    107738 to 107760 => 1860,
    107761 to 107782 => 1861,
    107783 to 107805 => 1862,
    107806 to 107827 => 1863,
    107828 to 107849 => 1864,
    107850 to 107872 => 1865,
    107873 to 107894 => 1866,
    107895 to 107916 => 1867,
    107917 to 107939 => 1868,
    107940 to 107961 => 1869,
    107962 to 107983 => 1870,
    107984 to 108005 => 1871,
    108006 to 108027 => 1872,
    108028 to 108050 => 1873,
    108051 to 108072 => 1874,
    108073 to 108094 => 1875,
    108095 to 108116 => 1876,
    108117 to 108138 => 1877,
    108139 to 108160 => 1878,
    108161 to 108182 => 1879,
    108183 to 108204 => 1880,
    108205 to 108226 => 1881,
    108227 to 108248 => 1882,
    108249 to 108270 => 1883,
    108271 to 108292 => 1884,
    108293 to 108314 => 1885,
    108315 to 108336 => 1886,
    108337 to 108358 => 1887,
    108359 to 108380 => 1888,
    108381 to 108402 => 1889,
    108403 to 108424 => 1890,
    108425 to 108446 => 1891,
    108447 to 108468 => 1892,
    108469 to 108489 => 1893,
    108490 to 108511 => 1894,
    108512 to 108533 => 1895,
    108534 to 108555 => 1896,
    108556 to 108577 => 1897,
    108578 to 108598 => 1898,
    108599 to 108620 => 1899,
    108621 to 108642 => 1900,
    108643 to 108663 => 1901,
    108664 to 108685 => 1902,
    108686 to 108707 => 1903,
    108708 to 108728 => 1904,
    108729 to 108750 => 1905,
    108751 to 108771 => 1906,
    108772 to 108793 => 1907,
    108794 to 108815 => 1908,
    108816 to 108836 => 1909,
    108837 to 108858 => 1910,
    108859 to 108879 => 1911,
    108880 to 108901 => 1912,
    108902 to 108922 => 1913,
    108923 to 108944 => 1914,
    108945 to 108965 => 1915,
    108966 to 108986 => 1916,
    108987 to 109008 => 1917,
    109009 to 109029 => 1918,
    109030 to 109050 => 1919,
    109051 to 109072 => 1920,
    109073 to 109093 => 1921,
    109094 to 109114 => 1922,
    109115 to 109136 => 1923,
    109137 to 109157 => 1924,
    109158 to 109178 => 1925,
    109179 to 109199 => 1926,
    109200 to 109221 => 1927,
    109222 to 109242 => 1928,
    109243 to 109263 => 1929,
    109264 to 109284 => 1930,
    109285 to 109305 => 1931,
    109306 to 109326 => 1932,
    109327 to 109348 => 1933,
    109349 to 109369 => 1934,
    109370 to 109390 => 1935,
    109391 to 109411 => 1936,
    109412 to 109432 => 1937,
    109433 to 109453 => 1938,
    109454 to 109474 => 1939,
    109475 to 109495 => 1940,
    109496 to 109516 => 1941,
    109517 to 109537 => 1942,
    109538 to 109558 => 1943,
    109559 to 109579 => 1944,
    109580 to 109600 => 1945,
    109601 to 109621 => 1946,
    109622 to 109641 => 1947,
    109642 to 109662 => 1948,
    109663 to 109683 => 1949,
    109684 to 109704 => 1950,
    109705 to 109725 => 1951,
    109726 to 109746 => 1952,
    109747 to 109766 => 1953,
    109767 to 109787 => 1954,
    109788 to 109808 => 1955,
    109809 to 109828 => 1956,
    109829 to 109849 => 1957,
    109850 to 109870 => 1958,
    109871 to 109891 => 1959,
    109892 to 109911 => 1960,
    109912 to 109932 => 1961,
    109933 to 109952 => 1962,
    109953 to 109973 => 1963,
    109974 to 109994 => 1964,
    109995 to 110014 => 1965,
    110015 to 110035 => 1966,
    110036 to 110055 => 1967,
    110056 to 110076 => 1968,
    110077 to 110096 => 1969,
    110097 to 110117 => 1970,
    110118 to 110137 => 1971,
    110138 to 110158 => 1972,
    110159 to 110178 => 1973,
    110179 to 110199 => 1974,
    110200 to 110219 => 1975,
    110220 to 110239 => 1976,
    110240 to 110260 => 1977,
    110261 to 110280 => 1978,
    110281 to 110300 => 1979,
    110301 to 110321 => 1980,
    110322 to 110341 => 1981,
    110342 to 110361 => 1982,
    110362 to 110382 => 1983,
    110383 to 110402 => 1984,
    110403 to 110422 => 1985,
    110423 to 110442 => 1986,
    110443 to 110463 => 1987,
    110464 to 110483 => 1988,
    110484 to 110503 => 1989,
    110504 to 110523 => 1990,
    110524 to 110543 => 1991,
    110544 to 110563 => 1992,
    110564 to 110584 => 1993,
    110585 to 110604 => 1994,
    110605 to 110624 => 1995,
    110625 to 110644 => 1996,
    110645 to 110664 => 1997,
    110665 to 110684 => 1998,
    110685 to 110704 => 1999,
    110705 to 110724 => 2000,
    110725 to 110744 => 2001,
    110745 to 110764 => 2002,
    110765 to 110784 => 2003,
    110785 to 110804 => 2004,
    110805 to 110824 => 2005,
    110825 to 110844 => 2006,
    110845 to 110863 => 2007,
    110864 to 110883 => 2008,
    110884 to 110903 => 2009,
    110904 to 110923 => 2010,
    110924 to 110943 => 2011,
    110944 to 110963 => 2012,
    110964 to 110982 => 2013,
    110983 to 111002 => 2014,
    111003 to 111022 => 2015,
    111023 to 111042 => 2016,
    111043 to 111061 => 2017,
    111062 to 111081 => 2018,
    111082 to 111101 => 2019,
    111102 to 111121 => 2020,
    111122 to 111140 => 2021,
    111141 to 111160 => 2022,
    111161 to 111179 => 2023,
    111180 to 111199 => 2024,
    111200 to 111219 => 2025,
    111220 to 111238 => 2026,
    111239 to 111258 => 2027,
    111259 to 111277 => 2028,
    111278 to 111297 => 2029,
    111298 to 111317 => 2030,
    111318 to 111336 => 2031,
    111337 to 111356 => 2032,
    111357 to 111375 => 2033,
    111376 to 111394 => 2034,
    111395 to 111414 => 2035,
    111415 to 111433 => 2036,
    111434 to 111453 => 2037,
    111454 to 111472 => 2038,
    111473 to 111492 => 2039,
    111493 to 111511 => 2040,
    111512 to 111530 => 2041,
    111531 to 111550 => 2042,
    111551 to 111569 => 2043,
    111570 to 111588 => 2044,
    111589 to 111608 => 2045,
    111609 to 111627 => 2046,
    111628 to 111637 => 2047
  );

 end package roi_atan;
