--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: Tube position coordinate
--  Multiplier: 32
--  Resolution: 0.03125 mm
--  
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TC_B_S3A_pkg is

  constant MAX_TUBES_INN : 5;
  constant MAX_TUBES_MID : 8;
  constant MAX_TUBES_OUT : 12;
  -- constant MAX_TUBES_EXT : 5;
  
  constant tube_coordinates_inn :  tube_coordinates_inn_aat(0 to MAX_TUBES_INN - 1)(0 to 7):= (
    --     layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       , layer 6       , layer 7       ,
    0 => ((      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100), -- tube 0
    1 => ((     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100), -- tube 1
    2 => ((    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100), -- tube 2
    3 => ((   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100), -- tube 3
    4 => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100)  -- tube 4
  );

  constant tube_coordinates_inn :  tube_coordinates_inn_aat(0 to MAX_TUBES_INN - 1)(0 to 6):= (
    --     layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       ,
    0 => ((      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100), -- tube 0
    1 => ((     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100), -- tube 1
    2 => ((    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100), -- tube 2
    3 => ((   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100), -- tube 3
    4 => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 4
    5 => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 5
    6 => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 6
    7 => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100)  -- tube 7
  );

  constant tube_coordinates_inn :  tube_coordinates_inn_aat(0 to MAX_TUBES_INN - 1)(0 to 6):= (
    --      layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       ,
    0  => ((      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100), -- tube 0
    1  => ((     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100), -- tube 1
    2  => ((    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100), -- tube 2
    3  => ((   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100), -- tube 3
    4  => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 4
    5  => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 5
    6  => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100), -- tube 6
    7  => ((  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100),(  10000,  100)  -- tube 7
    8  => ((      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100),(      1,  100), -- tube 8
    9  => ((     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100),(     10,  100), -- tube 9
    10 => ((    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100),(    100,  100), -- tube 10
    11 => ((   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100),(   1000,  100), -- tube 11

  );

  -- constant tube_coordinates_inn :  tube_coordinates_inn_aat(0 to MAX_TUBES_INN - 1)(0 to 7):= (

  -- );
  
  
end package TC_B_S3A_pkg;

