library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package board_pkg_common is

  --------------------------------------------------------------------------------
  -- MGT Mapping
  --------------------------------------------------------------------------------

  type gt_types_t is (GT_NIL, GTH, GTY);

  type mgt_types_t is (MGT_NIL, MGT_LPGBT_SIMPLEX, MGT_LPGBT, MGT_LPGBT_EMUL, MGT_C2C, MGT_SL, MGT_TCDS, MGT_FELIX);

  type mgt_inst_t is record
    mgt_type : mgt_types_t;
    refclk   : integer;
    gt_type  : gt_types_t;
    x_loc    : integer;
    y_loc    : integer;
  end record;

  type mgt_map_t is record
    mgt_id : integer;
  end record;

  type mgt_info_t is record
    gt_type      : gt_types_t;
    refclk0_freq : real;
    refclk1_freq : real;
  end record;

  constant c_mgtinfo_nil : mgt_info_t := (GT_NIL, 0.0, 0.0);
  constant c_mgt_nil     : mgt_inst_t := (MGT_NIL, -1, GT_NIL, -1, -1);

  type mgt_inst_array_t is array (integer range <>) of mgt_inst_t;
  type mgt_info_array_t is array (integer range <>) of mgt_info_t;
  type mgt_map_array_t is array (integer range <>) of mgt_map_t;

  --------------------------------------------------------------------------------
  -- REFCLK Mapping
  --------------------------------------------------------------------------------

  type refclk_types_t is (REFCLK_SYNC320, REFCLK_SYNC240, REFCLK_NIL);

  type refclk_types_array_t is array (integer range <>) of refclk_types_t;

  type station_id_t is (INNER, MIDDLE, OUTER, EXTRA);

  --------------------------------------------------------------------------------
  -- CSM Mapping
  --------------------------------------------------------------------------------

  type tdc_link_map_t is record
    link_id    : integer;
    elink      : integer;
    --enc_elink  : integer;
    station_id : integer;
    polmux_id  : integer;
    legacy     : boolean;
  end record;
  type tdc_link_map_array_t is array (integer range <>) of tdc_link_map_t;

  --------------------------------------------------------------------------------
  -- Utility Functions
  --------------------------------------------------------------------------------

  type int_array_t is array (integer range <>) of integer;

  function func_fill_subtype_idx (cnt_max : integer; mgt_list : mgt_inst_array_t; i_mgt_type : mgt_types_t; i_mgt_type_alt : mgt_types_t)
    return int_array_t;

  function func_count_link_types (mgt_list : mgt_inst_array_t; i_mgt_type : mgt_types_t)
    return integer;

  function func_count_tdc_links (tdc_map : tdc_link_map_array_t; mgt_list : mgt_inst_array_t)
    return integer;

  function func_count_polmux (tdc_map : tdc_link_map_array_t; num_tdcs : integer)
    return integer;

  function func_count_lpgbt_link_mapped_to_csm (tdc_map : tdc_link_map_array_t; num_tdcs : integer)
    return integer;

end package board_pkg_common;

package body board_pkg_common is

  function func_count_tdc_links (tdc_map : tdc_link_map_array_t; mgt_list : mgt_inst_array_t)
    return integer is
    variable count : integer := 0;
  begin
    for I in 0 to tdc_map'length-1 loop
      if (tdc_map(I).link_id >= 0) then
        assert ((mgt_list(tdc_map(I).link_id).mgt_type = MGT_LPGBT) or mgt_list(tdc_map(I).link_id).mgt_type = MGT_LPGBT_SIMPLEX) report "c_TDC_LINK_MAP specifies a tdc input on a non-lpgbt link" severity error;
        count := count + 1;
      end if;
    end loop;
    return count;
  end func_count_tdc_links;

  function func_fill_subtype_idx (cnt_max : integer; mgt_list : mgt_inst_array_t; i_mgt_type : mgt_types_t; i_mgt_type_alt : mgt_types_t)
    return int_array_t is
    variable count : integer := 0;
    variable idx   : int_array_t (0 to mgt_list'length-1);
  begin
    for I in 0 to mgt_list'length-1 loop
      if (count < cnt_max and (mgt_list(I).mgt_type = i_mgt_type or mgt_list(I).mgt_type = i_mgt_type_alt)) then
        idx(I) := count;
        count  := count + 1;
      else
        idx(I) := -1;
      end if;
    end loop;  -- I
    return idx;
  end func_fill_subtype_idx;

  function func_count_link_types (mgt_list : mgt_inst_array_t; i_mgt_type : mgt_types_t)
    return integer is
    variable count : integer := 0;
  begin
    for I in 0 to mgt_list'length-1 loop
      if (mgt_list(I).mgt_type = i_mgt_type) then
        count := count + 1;
      end if;
    end loop;
    return count;
  end func_count_link_types;

  -- write function to count number of polmuxes
  function func_count_polmux (tdc_map : tdc_link_map_array_t; num_tdcs : integer)
    return integer is
    variable max : integer := 0;
  begin
    for I in 0 to num_tdcs-1 loop
      if (tdc_map(I).polmux_id > max) then
        max := tdc_map(I).polmux_id;
      end if;
    end loop;
    return max+1; -- the count is the index of the highest number + 1
  end func_count_polmux;

  -- write function to count number of polmuxes
  function func_count_lpgbt_link_mapped_to_csm (tdc_map : tdc_link_map_array_t; num_tdcs : integer)
    return integer is
    variable max : integer := 0;
  begin
    for I in 0 to num_tdcs-1 loop
      if (tdc_map(I).link_id > max) then
        max := tdc_map(I).link_id;
      end if;
    end loop;
    return max+1;
  end func_count_lpgbt_link_mapped_to_csm;

end package body;
