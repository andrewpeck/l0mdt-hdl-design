library ieee;
use ieee.std_logic_1164.all;

package fullmode_pkg is

  type std_logic_vector_array is array(integer range <>) of std_logic_vector;
  
end package fullmode_pkg;
