--------------------------------------------------------------------------------
-- UMass , Physics Department
-- Project: ATLAS L0MDT Trigger
-- File: apb_pkg.vhd
-- Module: <<moduleName>>
-- File PATH: /shared/APBus/pkg/apb_pkg.vhd
-- -----
-- File Created: Monday, 12th July 2021 12:20:43 pm
-- Author: Guillermo Loustau de Linares (guillermo.ldl@cern.ch)
-- -----
-- Last Modified: Thursday, 16th December 2021 12:06:22 am
-- Modified By: Guillermo Loustau de Linares (guillermo.ldl@cern.ch>)
-- -----
-- HISTORY:
--------------------------------------------------------------------------------



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package apb_pkg is
  
  constant c_DUMMY : integer := 0;
  
  
end package apb_pkg;

package body apb_pkg is
  
  
  
  
end package body apb_pkg;
