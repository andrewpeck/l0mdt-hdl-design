library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;
use std.standard.all;
use std.textio.all;

package pt_params_pkg is
-- ComboId to ROM index function declaration
function comboid_to_index_ram(comboid : unsigned) return std_logic_vector;

-- pT parametrisation constants
constant params_width : natural := 32;
constant a0_width     : natural := 11;
constant a1_width     : natural := 23;
constant b0_width     : natural := 12;
constant b1_width     : natural := 8;
constant b2_width     : natural := 4;
constant c0_width     : natural := 16;
constant c1_width     : natural := 6;

constant params_depth_width : natural := 9;
 
type t_params is
record 
    a0              :  signed(params_width-1 downto 0);
    a1              :  signed(params_width-1 downto 0);
    b0              :  signed(params_width-1 downto 0);
    b1              :  signed(params_width-1 downto 0);
    b2              :  signed(params_width-1 downto 0);
    c0              :  signed(params_width-1 downto 0);
    c1              :  signed(params_width-1 downto 0);
end record;

constant null_params : t_params    := ((others => '0') , (others => '0'), (others => '0'), (others => '0'), (others => '0'), (others => '0'), (others => '0'));
--RAM containing pT parametrisation constants

type t_params_ram is array(511 downto 0) of t_params;
function pt_parameter return t_params_ram;
end;
package body pt_params_pkg is

-- ComboId to ROM index function body
function comboid_to_index_ram(comboid : unsigned) return std_logic_vector is
   variable index : integer := 0;
   variable addr : std_logic_vector(params_depth_width-1 downto 0);
begin
   if comboid = 10 then
       index := 0;
   end if;
   if comboid = 522 then
       index := 1;
   end if;
   if comboid = 1034 then
       index := 2;
   end if;
   if comboid = 1546 then
       index := 3;
   end if;
   if comboid = 2058 then
       index := 4;
   end if;
   if comboid = 2570 then
       index := 5;
   end if;
   if comboid = 3082 then
       index := 6;
   end if;
   if comboid = 3594 then
       index := 7;
   end if;
   if comboid = 4106 then
       index := 8;
   end if;
   if comboid = 4618 then
       index := 9;
   end if;
   if comboid = 130 then
       index := 10;
   end if;
   if comboid = 642 then
       index := 11;
   end if;
   if comboid = 1154 then
       index := 12;
   end if;
   if comboid = 1666 then
       index := 13;
   end if;
   if comboid = 2178 then
       index := 14;
   end if;
   if comboid = 2690 then
       index := 15;
   end if;
   if comboid = 3202 then
       index := 16;
   end if;
   if comboid = 3714 then
       index := 17;
   end if;
   if comboid = 4226 then
       index := 18;
   end if;
   if comboid = 4738 then
       index := 19;
   end if;
   if comboid = 138 then
       index := 20;
   end if;
   if comboid = 650 then
       index := 21;
   end if;
   if comboid = 1162 then
       index := 22;
   end if;
   if comboid = 1674 then
       index := 23;
   end if;
   if comboid = 2186 then
       index := 24;
   end if;
   if comboid = 2698 then
       index := 25;
   end if;
   if comboid = 3210 then
       index := 26;
   end if;
   if comboid = 3722 then
       index := 27;
   end if;
   if comboid = 4234 then
       index := 28;
   end if;
   if comboid = 4746 then
       index := 29;
   end if;
   if comboid = 146 then
       index := 30;
   end if;
   if comboid = 658 then
       index := 31;
   end if;
   if comboid = 1170 then
       index := 32;
   end if;
   if comboid = 1682 then
       index := 33;
   end if;
   if comboid = 2194 then
       index := 34;
   end if;
   if comboid = 2706 then
       index := 35;
   end if;
   if comboid = 3218 then
       index := 36;
   end if;
   if comboid = 3730 then
       index := 37;
   end if;
   if comboid = 4242 then
       index := 38;
   end if;
   if comboid = 4754 then
       index := 39;
   end if;
   if comboid = 147 then
       index := 40;
   end if;
   if comboid = 659 then
       index := 41;
   end if;
   if comboid = 1171 then
       index := 42;
   end if;
   if comboid = 1683 then
       index := 43;
   end if;
   if comboid = 2195 then
       index := 44;
   end if;
   if comboid = 2707 then
       index := 45;
   end if;
   if comboid = 3219 then
       index := 46;
   end if;
   if comboid = 3731 then
       index := 47;
   end if;
   if comboid = 4243 then
       index := 48;
   end if;
   if comboid = 4755 then
       index := 49;
   end if;
   if comboid = 18 then
       index := 50;
   end if;
   if comboid = 530 then
       index := 51;
   end if;
   if comboid = 1042 then
       index := 52;
   end if;
   if comboid = 1554 then
       index := 53;
   end if;
   if comboid = 2066 then
       index := 54;
   end if;
   if comboid = 2578 then
       index := 55;
   end if;
   if comboid = 3090 then
       index := 56;
   end if;
   if comboid = 3602 then
       index := 57;
   end if;
   if comboid = 4114 then
       index := 58;
   end if;
   if comboid = 4626 then
       index := 59;
   end if;
   if comboid = 19 then
       index := 60;
   end if;
   if comboid = 531 then
       index := 61;
   end if;
   if comboid = 1043 then
       index := 62;
   end if;
   if comboid = 1555 then
       index := 63;
   end if;
   if comboid = 2067 then
       index := 64;
   end if;
   if comboid = 2579 then
       index := 65;
   end if;
   if comboid = 3091 then
       index := 66;
   end if;
   if comboid = 3603 then
       index := 67;
   end if;
   if comboid = 4115 then
       index := 68;
   end if;
   if comboid = 4627 then
       index := 69;
   end if;
   if comboid = 195 then
       index := 70;
   end if;
   if comboid = 707 then
       index := 71;
   end if;
   if comboid = 1219 then
       index := 72;
   end if;
   if comboid = 1731 then
       index := 73;
   end if;
   if comboid = 2243 then
       index := 74;
   end if;
   if comboid = 2755 then
       index := 75;
   end if;
   if comboid = 3267 then
       index := 76;
   end if;
   if comboid = 3779 then
       index := 77;
   end if;
   if comboid = 4291 then
       index := 78;
   end if;
   if comboid = 4803 then
       index := 79;
   end if;
   if comboid = 210 then
       index := 80;
   end if;
   if comboid = 722 then
       index := 81;
   end if;
   if comboid = 1234 then
       index := 82;
   end if;
   if comboid = 1746 then
       index := 83;
   end if;
   if comboid = 2258 then
       index := 84;
   end if;
   if comboid = 2770 then
       index := 85;
   end if;
   if comboid = 3282 then
       index := 86;
   end if;
   if comboid = 3794 then
       index := 87;
   end if;
   if comboid = 4306 then
       index := 88;
   end if;
   if comboid = 4818 then
       index := 89;
   end if;
   if comboid = 211 then
       index := 90;
   end if;
   if comboid = 723 then
       index := 91;
   end if;
   if comboid = 1235 then
       index := 92;
   end if;
   if comboid = 1747 then
       index := 93;
   end if;
   if comboid = 2259 then
       index := 94;
   end if;
   if comboid = 2771 then
       index := 95;
   end if;
   if comboid = 3283 then
       index := 96;
   end if;
   if comboid = 3795 then
       index := 97;
   end if;
   if comboid = 4307 then
       index := 98;
   end if;
   if comboid = 4819 then
       index := 99;
   end if;
   if comboid = 219 then
       index := 100;
   end if;
   if comboid = 731 then
       index := 101;
   end if;
   if comboid = 1243 then
       index := 102;
   end if;
   if comboid = 1755 then
       index := 103;
   end if;
   if comboid = 2267 then
       index := 104;
   end if;
   if comboid = 2779 then
       index := 105;
   end if;
   if comboid = 3291 then
       index := 106;
   end if;
   if comboid = 3803 then
       index := 107;
   end if;
   if comboid = 4315 then
       index := 108;
   end if;
   if comboid = 4827 then
       index := 109;
   end if;
   if comboid = 27 then
       index := 110;
   end if;
   if comboid = 539 then
       index := 111;
   end if;
   if comboid = 1051 then
       index := 112;
   end if;
   if comboid = 1563 then
       index := 113;
   end if;
   if comboid = 2075 then
       index := 114;
   end if;
   if comboid = 2587 then
       index := 115;
   end if;
   if comboid = 3099 then
       index := 116;
   end if;
   if comboid = 3611 then
       index := 117;
   end if;
   if comboid = 4123 then
       index := 118;
   end if;
   if comboid = 4635 then
       index := 119;
   end if;
   if comboid = 28 then
       index := 120;
   end if;
   if comboid = 540 then
       index := 121;
   end if;
   if comboid = 1052 then
       index := 122;
   end if;
   if comboid = 1564 then
       index := 123;
   end if;
   if comboid = 2076 then
       index := 124;
   end if;
   if comboid = 2588 then
       index := 125;
   end if;
   if comboid = 3100 then
       index := 126;
   end if;
   if comboid = 3612 then
       index := 127;
   end if;
   if comboid = 4124 then
       index := 128;
   end if;
   if comboid = 4636 then
       index := 129;
   end if;
   if comboid = 280 then
       index := 130;
   end if;
   if comboid = 792 then
       index := 131;
   end if;
   if comboid = 1304 then
       index := 132;
   end if;
   if comboid = 1816 then
       index := 133;
   end if;
   if comboid = 2328 then
       index := 134;
   end if;
   if comboid = 2840 then
       index := 135;
   end if;
   if comboid = 3352 then
       index := 136;
   end if;
   if comboid = 3864 then
       index := 137;
   end if;
   if comboid = 4376 then
       index := 138;
   end if;
   if comboid = 4888 then
       index := 139;
   end if;
   if comboid = 283 then
       index := 140;
   end if;
   if comboid = 795 then
       index := 141;
   end if;
   if comboid = 1307 then
       index := 142;
   end if;
   if comboid = 1819 then
       index := 143;
   end if;
   if comboid = 2331 then
       index := 144;
   end if;
   if comboid = 2843 then
       index := 145;
   end if;
   if comboid = 3355 then
       index := 146;
   end if;
   if comboid = 3867 then
       index := 147;
   end if;
   if comboid = 4379 then
       index := 148;
   end if;
   if comboid = 4891 then
       index := 149;
   end if;
   if comboid = 284 then
       index := 150;
   end if;
   if comboid = 796 then
       index := 151;
   end if;
   if comboid = 1308 then
       index := 152;
   end if;
   if comboid = 1820 then
       index := 153;
   end if;
   if comboid = 2332 then
       index := 154;
   end if;
   if comboid = 2844 then
       index := 155;
   end if;
   if comboid = 3356 then
       index := 156;
   end if;
   if comboid = 3868 then
       index := 157;
   end if;
   if comboid = 4380 then
       index := 158;
   end if;
   if comboid = 4892 then
       index := 159;
   end if;
   if comboid = 292 then
       index := 160;
   end if;
   if comboid = 804 then
       index := 161;
   end if;
   if comboid = 1316 then
       index := 162;
   end if;
   if comboid = 1828 then
       index := 163;
   end if;
   if comboid = 2340 then
       index := 164;
   end if;
   if comboid = 2852 then
       index := 165;
   end if;
   if comboid = 3364 then
       index := 166;
   end if;
   if comboid = 3876 then
       index := 167;
   end if;
   if comboid = 4388 then
       index := 168;
   end if;
   if comboid = 4900 then
       index := 169;
   end if;
   if comboid = 356 then
       index := 170;
   end if;
   if comboid = 868 then
       index := 171;
   end if;
   if comboid = 1380 then
       index := 172;
   end if;
   if comboid = 1892 then
       index := 173;
   end if;
   if comboid = 2404 then
       index := 174;
   end if;
   if comboid = 2916 then
       index := 175;
   end if;
   if comboid = 3428 then
       index := 176;
   end if;
   if comboid = 3940 then
       index := 177;
   end if;
   if comboid = 4452 then
       index := 178;
   end if;
   if comboid = 4964 then
       index := 179;
   end if;
   if comboid = 36 then
       index := 180;
   end if;
   if comboid = 548 then
       index := 181;
   end if;
   if comboid = 1060 then
       index := 182;
   end if;
   if comboid = 1572 then
       index := 183;
   end if;
   if comboid = 2084 then
       index := 184;
   end if;
   if comboid = 2596 then
       index := 185;
   end if;
   if comboid = 3108 then
       index := 186;
   end if;
   if comboid = 3620 then
       index := 187;
   end if;
   if comboid = 4132 then
       index := 188;
   end if;
   if comboid = 4644 then
       index := 189;
   end if;
   if comboid = 364 then
       index := 190;
   end if;
   if comboid = 876 then
       index := 191;
   end if;
   if comboid = 1388 then
       index := 192;
   end if;
   if comboid = 1900 then
       index := 193;
   end if;
   if comboid = 2412 then
       index := 194;
   end if;
   if comboid = 2924 then
       index := 195;
   end if;
   if comboid = 3436 then
       index := 196;
   end if;
   if comboid = 3948 then
       index := 197;
   end if;
   if comboid = 4460 then
       index := 198;
   end if;
   if comboid = 4972 then
       index := 199;
   end if;
   if comboid = 365 then
       index := 200;
   end if;
   if comboid = 877 then
       index := 201;
   end if;
   if comboid = 1389 then
       index := 202;
   end if;
   if comboid = 1901 then
       index := 203;
   end if;
   if comboid = 2413 then
       index := 204;
   end if;
   if comboid = 2925 then
       index := 205;
   end if;
   if comboid = 3437 then
       index := 206;
   end if;
   if comboid = 3949 then
       index := 207;
   end if;
   if comboid = 4461 then
       index := 208;
   end if;
   if comboid = 4973 then
       index := 209;
   end if;
   if comboid = 373 then
       index := 210;
   end if;
   if comboid = 885 then
       index := 211;
   end if;
   if comboid = 1397 then
       index := 212;
   end if;
   if comboid = 1909 then
       index := 213;
   end if;
   if comboid = 2421 then
       index := 214;
   end if;
   if comboid = 2933 then
       index := 215;
   end if;
   if comboid = 3445 then
       index := 216;
   end if;
   if comboid = 3957 then
       index := 217;
   end if;
   if comboid = 4469 then
       index := 218;
   end if;
   if comboid = 4981 then
       index := 219;
   end if;
   if comboid = 374 then
       index := 220;
   end if;
   if comboid = 886 then
       index := 221;
   end if;
   if comboid = 1398 then
       index := 222;
   end if;
   if comboid = 1910 then
       index := 223;
   end if;
   if comboid = 2422 then
       index := 224;
   end if;
   if comboid = 2934 then
       index := 225;
   end if;
   if comboid = 3446 then
       index := 226;
   end if;
   if comboid = 3958 then
       index := 227;
   end if;
   if comboid = 4470 then
       index := 228;
   end if;
   if comboid = 4982 then
       index := 229;
   end if;
   if comboid = 390 then
       index := 230;
   end if;
   if comboid = 902 then
       index := 231;
   end if;
   if comboid = 1414 then
       index := 232;
   end if;
   if comboid = 1926 then
       index := 233;
   end if;
   if comboid = 2438 then
       index := 234;
   end if;
   if comboid = 2950 then
       index := 235;
   end if;
   if comboid = 3462 then
       index := 236;
   end if;
   if comboid = 3974 then
       index := 237;
   end if;
   if comboid = 4486 then
       index := 238;
   end if;
   if comboid = 4998 then
       index := 239;
   end if;
   if comboid = 438 then
       index := 240;
   end if;
   if comboid = 950 then
       index := 241;
   end if;
   if comboid = 1462 then
       index := 242;
   end if;
   if comboid = 1974 then
       index := 243;
   end if;
   if comboid = 2486 then
       index := 244;
   end if;
   if comboid = 2998 then
       index := 245;
   end if;
   if comboid = 3510 then
       index := 246;
   end if;
   if comboid = 4022 then
       index := 247;
   end if;
   if comboid = 4534 then
       index := 248;
   end if;
   if comboid = 5046 then
       index := 249;
   end if;
   if comboid = 45 then
       index := 250;
   end if;
   if comboid = 557 then
       index := 251;
   end if;
   if comboid = 1069 then
       index := 252;
   end if;
   if comboid = 1581 then
       index := 253;
   end if;
   if comboid = 2093 then
       index := 254;
   end if;
   if comboid = 2605 then
       index := 255;
   end if;
   if comboid = 3117 then
       index := 256;
   end if;
   if comboid = 3629 then
       index := 257;
   end if;
   if comboid = 4141 then
       index := 258;
   end if;
   if comboid = 4653 then
       index := 259;
   end if;
   if comboid = 53 then
       index := 260;
   end if;
   if comboid = 565 then
       index := 261;
   end if;
   if comboid = 1077 then
       index := 262;
   end if;
   if comboid = 1589 then
       index := 263;
   end if;
   if comboid = 2101 then
       index := 264;
   end if;
   if comboid = 2613 then
       index := 265;
   end if;
   if comboid = 3125 then
       index := 266;
   end if;
   if comboid = 3637 then
       index := 267;
   end if;
   if comboid = 4149 then
       index := 268;
   end if;
   if comboid = 4661 then
       index := 269;
   end if;
   if comboid = 54 then
       index := 270;
   end if;
   if comboid = 566 then
       index := 271;
   end if;
   if comboid = 1078 then
       index := 272;
   end if;
   if comboid = 1590 then
       index := 273;
   end if;
   if comboid = 2102 then
       index := 274;
   end if;
   if comboid = 2614 then
       index := 275;
   end if;
   if comboid = 3126 then
       index := 276;
   end if;
   if comboid = 3638 then
       index := 277;
   end if;
   if comboid = 4150 then
       index := 278;
   end if;
   if comboid = 4662 then
       index := 279;
   end if;
   if comboid = 66 then
       index := 280;
   end if;
   if comboid = 578 then
       index := 281;
   end if;
   if comboid = 1090 then
       index := 282;
   end if;
   if comboid = 1602 then
       index := 283;
   end if;
   if comboid = 2114 then
       index := 284;
   end if;
   if comboid = 2626 then
       index := 285;
   end if;
   if comboid = 3138 then
       index := 286;
   end if;
   if comboid = 3650 then
       index := 287;
   end if;
   if comboid = 4162 then
       index := 288;
   end if;
   if comboid = 4674 then
       index := 289;
   end if;
   if comboid = 72 then
       index := 290;
   end if;
   if comboid = 584 then
       index := 291;
   end if;
   if comboid = 1096 then
       index := 292;
   end if;
   if comboid = 1608 then
       index := 293;
   end if;
   if comboid = 2120 then
       index := 294;
   end if;
   if comboid = 2632 then
       index := 295;
   end if;
   if comboid = 3144 then
       index := 296;
   end if;
   if comboid = 3656 then
       index := 297;
   end if;
   if comboid = 4168 then
       index := 298;
   end if;
   if comboid = 4680 then
       index := 299;
   end if;
   if comboid = 74 then
       index := 300;
   end if;
   if comboid = 586 then
       index := 301;
   end if;
   if comboid = 1098 then
       index := 302;
   end if;
   if comboid = 1610 then
       index := 303;
   end if;
   if comboid = 2122 then
       index := 304;
   end if;
   if comboid = 2634 then
       index := 305;
   end if;
   if comboid = 3146 then
       index := 306;
   end if;
   if comboid = 3658 then
       index := 307;
   end if;
   if comboid = 4170 then
       index := 308;
   end if;
   if comboid = 4682 then
       index := 309;
   end if;
   
   addr := std_logic_vector(to_unsigned(index, params_depth_width));
   return addr;
end function;

function pt_parameter return t_params_ram is 
   variable ram : t_params_ram := (others => null_params);
begin
   ram(0) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(1) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(75, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(10, params_width), to_signed(0, params_width));
   ram(2) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(125, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(7, params_width), to_signed(0, params_width));
   ram(3) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(135, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(26, params_width), to_signed(0, params_width));
   ram(4) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(186, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(69, params_width), to_signed(0, params_width));
   ram(5) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(278, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-53, params_width), to_signed(0, params_width));
   ram(6) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(298, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(49, params_width), to_signed(0, params_width));
   ram(7) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(405, params_width), to_signed(3, params_width), to_signed(-2, params_width), to_signed(-62, params_width), to_signed(0, params_width));
   ram(8) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(394, params_width), to_signed(5, params_width), to_signed(-2, params_width), to_signed(-165, params_width), to_signed(0, params_width));
   ram(9) := ( to_signed(309, params_width), to_signed(2131, params_width), to_signed(618, params_width), to_signed(3, params_width), to_signed(0, params_width), to_signed(96, params_width), to_signed(1, params_width));
   ram(10) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(11) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(174, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(71, params_width), to_signed(0, params_width));
   ram(12) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(198, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(46, params_width), to_signed(0, params_width));
   ram(13) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(181, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(145, params_width), to_signed(0, params_width));
   ram(14) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(222, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(89, params_width), to_signed(0, params_width));
   ram(15) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(135, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-63, params_width), to_signed(0, params_width));
   ram(16) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(129, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(79, params_width), to_signed(0, params_width));
   ram(17) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(263, params_width), to_signed(2, params_width), to_signed(-1, params_width), to_signed(51, params_width), to_signed(0, params_width));
   ram(18) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(245, params_width), to_signed(-3, params_width), to_signed(-2, params_width), to_signed(80, params_width), to_signed(0, params_width));
   ram(19) := ( to_signed(430, params_width), to_signed(3592, params_width), to_signed(201, params_width), to_signed(5, params_width), to_signed(-1, params_width), to_signed(320, params_width), to_signed(-1, params_width));
   ram(20) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(21) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(134, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(260, params_width), to_signed(-1, params_width));
   ram(22) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(84, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(438, params_width), to_signed(-1, params_width));
   ram(23) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(98, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(161, params_width), to_signed(0, params_width));
   ram(24) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(155, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-165, params_width), to_signed(0, params_width));
   ram(25) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(133, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(375, params_width), to_signed(-1, params_width));
   ram(26) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(142, params_width), to_signed(-5, params_width), to_signed(-1, params_width), to_signed(-191, params_width), to_signed(0, params_width));
   ram(27) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(10, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(-482, params_width), to_signed(1, params_width));
   ram(28) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(147, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(-975, params_width), to_signed(2, params_width));
   ram(29) := ( to_signed(384, params_width), to_signed(2257856, params_width), to_signed(273, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-112, params_width), to_signed(0, params_width));
   ram(30) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(31) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(128, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-20, params_width), to_signed(0, params_width));
   ram(32) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(132, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(87, params_width), to_signed(0, params_width));
   ram(33) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(129, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(101, params_width), to_signed(0, params_width));
   ram(34) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(140, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(185, params_width), to_signed(0, params_width));
   ram(35) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(143, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(286, params_width), to_signed(0, params_width));
   ram(36) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(146, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(338, params_width), to_signed(-1, params_width));
   ram(37) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(156, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(405, params_width), to_signed(-1, params_width));
   ram(38) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(145, params_width), to_signed(-1, params_width), to_signed(-2, params_width), to_signed(400, params_width), to_signed(-1, params_width));
   ram(39) := ( to_signed(403, params_width), to_signed(2332320, params_width), to_signed(249, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(439, params_width), to_signed(-1, params_width));
   ram(40) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(41) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(80, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(84, params_width), to_signed(0, params_width));
   ram(42) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(87, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(328, params_width), to_signed(0, params_width));
   ram(43) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(95, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-972, params_width), to_signed(1, params_width));
   ram(44) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(174, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-988, params_width), to_signed(1, params_width));
   ram(45) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(46) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(47) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(48) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(49) := ( to_signed(302, params_width), to_signed(2492621, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(50) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(51) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(95, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-52, params_width), to_signed(0, params_width));
   ram(52) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(124, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(22, params_width), to_signed(0, params_width));
   ram(53) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(169, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-9, params_width), to_signed(0, params_width));
   ram(54) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(237, params_width), to_signed(-6, params_width), to_signed(-1, params_width), to_signed(310, params_width), to_signed(0, params_width));
   ram(55) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(277, params_width), to_signed(-8, params_width), to_signed(-2, params_width), to_signed(518, params_width), to_signed(-1, params_width));
   ram(56) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(296, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(524, params_width), to_signed(-1, params_width));
   ram(57) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(319, params_width), to_signed(12, params_width), to_signed(0, params_width), to_signed(507, params_width), to_signed(-1, params_width));
   ram(58) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(541, params_width), to_signed(10, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(59) := ( to_signed(325, params_width), to_signed(2136, params_width), to_signed(939, params_width), to_signed(19, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(60) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(61) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(58, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(203, params_width), to_signed(0, params_width));
   ram(62) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(158, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(-2416, params_width), to_signed(3, params_width));
   ram(63) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(245, params_width), to_signed(4, params_width), to_signed(-1, params_width), to_signed(5543, params_width), to_signed(-7, params_width));
   ram(64) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(287, params_width), to_signed(-2, params_width), to_signed(-2, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(65) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(66) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(350, params_width), to_signed(10, params_width), to_signed(-4, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(67) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(68) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(69) := ( to_signed(339, params_width), to_signed(2086, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(70) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(71) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(141, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-159, params_width), to_signed(0, params_width));
   ram(72) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(152, params_width), to_signed(2, params_width), to_signed(-1, params_width), to_signed(-222, params_width), to_signed(0, params_width));
   ram(73) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(195, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(-338, params_width), to_signed(0, params_width));
   ram(74) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(164, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(61, params_width), to_signed(0, params_width));
   ram(75) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(142, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-95, params_width), to_signed(0, params_width));
   ram(76) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(271, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-790, params_width), to_signed(1, params_width));
   ram(77) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(204, params_width), to_signed(7, params_width), to_signed(-1, params_width), to_signed(848, params_width), to_signed(-1, params_width));
   ram(78) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(372, params_width), to_signed(3, params_width), to_signed(-2, params_width), to_signed(-284, params_width), to_signed(0, params_width));
   ram(79) := ( to_signed(391, params_width), to_signed(3641, params_width), to_signed(357, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(-182, params_width), to_signed(0, params_width));
   ram(80) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(81) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(110, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(978, params_width), to_signed(-1, params_width));
   ram(82) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(103, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(340, params_width), to_signed(0, params_width));
   ram(83) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(101, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(1010, params_width), to_signed(-1, params_width));
   ram(84) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(143, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(1905, params_width), to_signed(-3, params_width));
   ram(85) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(113, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(-3908, params_width), to_signed(5, params_width));
   ram(86) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(-86, params_width), to_signed(3, params_width), to_signed(-1, params_width), to_signed(3112, params_width), to_signed(-4, params_width));
   ram(87) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(54, params_width), to_signed(-4, params_width), to_signed(-2, params_width), to_signed(-328, params_width), to_signed(0, params_width));
   ram(88) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(40, params_width), to_signed(-6, params_width), to_signed(-1, params_width), to_signed(-1278, params_width), to_signed(2, params_width));
   ram(89) := ( to_signed(432, params_width), to_signed(2327642, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(90) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(91) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(92) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(192, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(455, params_width), to_signed(-1, params_width));
   ram(93) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(118, params_width), to_signed(2, params_width), to_signed(-1, params_width), to_signed(-1320, params_width), to_signed(2, params_width));
   ram(94) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(50, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-1862, params_width), to_signed(2, params_width));
   ram(95) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(-43, params_width), to_signed(2, params_width), to_signed(-1, params_width), to_signed(-1252, params_width), to_signed(2, params_width));
   ram(96) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(-98, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(190, params_width), to_signed(0, params_width));
   ram(97) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(-181, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(30, params_width), to_signed(0, params_width));
   ram(98) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(-196, params_width), to_signed(-5, params_width), to_signed(-1, params_width), to_signed(403, params_width), to_signed(0, params_width));
   ram(99) := ( to_signed(610, params_width), to_signed(2057677, params_width), to_signed(-129, params_width), to_signed(3, params_width), to_signed(0, params_width), to_signed(512, params_width), to_signed(-1, params_width));
   ram(100) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(101) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(137, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-101, params_width), to_signed(0, params_width));
   ram(102) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(124, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(158, params_width), to_signed(0, params_width));
   ram(103) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(113, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(408, params_width), to_signed(0, params_width));
   ram(104) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(98, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(525, params_width), to_signed(-1, params_width));
   ram(105) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(116, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(898, params_width), to_signed(-1, params_width));
   ram(106) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(107, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(927, params_width), to_signed(-1, params_width));
   ram(107) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(106, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(1238, params_width), to_signed(-1, params_width));
   ram(108) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(124, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(1024, params_width), to_signed(-1, params_width));
   ram(109) := ( to_signed(415, params_width), to_signed(2493760, params_width), to_signed(245, params_width), to_signed(-5, params_width), to_signed(-1, params_width), to_signed(857, params_width), to_signed(-1, params_width));
   ram(110) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(111) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(88, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(109, params_width), to_signed(0, params_width));
   ram(112) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(148, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(5, params_width), to_signed(0, params_width));
   ram(113) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(190, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(214, params_width), to_signed(0, params_width));
   ram(114) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(227, params_width), to_signed(-7, params_width), to_signed(-1, params_width), to_signed(779, params_width), to_signed(-1, params_width));
   ram(115) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(354, params_width), to_signed(-2, params_width), to_signed(-2, params_width), to_signed(1209, params_width), to_signed(-1, params_width));
   ram(116) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(302, params_width), to_signed(-11, params_width), to_signed(0, params_width), to_signed(-194, params_width), to_signed(0, params_width));
   ram(117) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(125, params_width), to_signed(82, params_width), to_signed(2, params_width), to_signed(2154, params_width), to_signed(-2, params_width));
   ram(118) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(471, params_width), to_signed(24, params_width), to_signed(3, params_width), to_signed(-290, params_width), to_signed(1, params_width));
   ram(119) := ( to_signed(351, params_width), to_signed(2152, params_width), to_signed(1733, params_width), to_signed(34, params_width), to_signed(-2, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(120) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(121) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(80, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(-667, params_width), to_signed(1, params_width));
   ram(122) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(19, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-1588, params_width), to_signed(1, params_width));
   ram(123) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(98, params_width), to_signed(-9, params_width), to_signed(-2, params_width), to_signed(-569, params_width), to_signed(1, params_width));
   ram(124) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(180, params_width), to_signed(17, params_width), to_signed(-1, params_width), to_signed(909, params_width), to_signed(-1, params_width));
   ram(125) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(183, params_width), to_signed(38, params_width), to_signed(1, params_width), to_signed(3941, params_width), to_signed(-4, params_width));
   ram(126) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-9813, params_width), to_signed(9, params_width));
   ram(127) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(128) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(129) := ( to_signed(326, params_width), to_signed(1967, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(130) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(131) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(132) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(309, params_width), to_signed(-21, params_width), to_signed(-2, params_width), to_signed(-1556, params_width), to_signed(1, params_width));
   ram(133) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(468, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(-2068, params_width), to_signed(2, params_width));
   ram(134) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(518, params_width), to_signed(-7, params_width), to_signed(-2, params_width), to_signed(-440, params_width), to_signed(0, params_width));
   ram(135) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(592, params_width), to_signed(-11, params_width), to_signed(-3, params_width), to_signed(-3456, params_width), to_signed(3, params_width));
   ram(136) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(567, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(-182, params_width), to_signed(0, params_width));
   ram(137) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(656, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(1350, params_width), to_signed(-1, params_width));
   ram(138) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(701, params_width), to_signed(5, params_width), to_signed(-1, params_width), to_signed(-368, params_width), to_signed(0, params_width));
   ram(139) := ( to_signed(650, params_width), to_signed(1786, params_width), to_signed(928, params_width), to_signed(3, params_width), to_signed(0, params_width), to_signed(-277, params_width), to_signed(1, params_width));
   ram(140) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(141) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(180, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(335, params_width), to_signed(0, params_width));
   ram(142) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(145, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-75, params_width), to_signed(0, params_width));
   ram(143) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(91, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-251, params_width), to_signed(0, params_width));
   ram(144) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(85, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-2064, params_width), to_signed(2, params_width));
   ram(145) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(45, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-5393, params_width), to_signed(5, params_width));
   ram(146) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(20, params_width), to_signed(-1, params_width), to_signed(-2, params_width), to_signed(-6772, params_width), to_signed(6, params_width));
   ram(147) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(-37, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(-7114, params_width), to_signed(7, params_width));
   ram(148) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(-111, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-5948, params_width), to_signed(5, params_width));
   ram(149) := ( to_signed(519, params_width), to_signed(2427731, params_width), to_signed(133, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-6771, params_width), to_signed(6, params_width));
   ram(150) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(151) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(81, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-1762, params_width), to_signed(2, params_width));
   ram(152) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(103, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(984, params_width), to_signed(-1, params_width));
   ram(153) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(100, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(1588, params_width), to_signed(-1, params_width));
   ram(154) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(91, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(3606, params_width), to_signed(-3, params_width));
   ram(155) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(91, params_width), to_signed(3, params_width), to_signed(-1, params_width), to_signed(4262, params_width), to_signed(-4, params_width));
   ram(156) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(82, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(6679, params_width), to_signed(-6, params_width));
   ram(157) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(67, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(4357, params_width), to_signed(-4, params_width));
   ram(158) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(74, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(7229, params_width), to_signed(-6, params_width));
   ram(159) := ( to_signed(397, params_width), to_signed(2528486, params_width), to_signed(120, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(6968, params_width), to_signed(-6, params_width));
   ram(160) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(161) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(153, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(-458, params_width), to_signed(0, params_width));
   ram(162) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(135, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-331, params_width), to_signed(0, params_width));
   ram(163) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(105, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(70, params_width), to_signed(0, params_width));
   ram(164) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(96, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(410, params_width), to_signed(0, params_width));
   ram(165) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(76, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(725, params_width), to_signed(-1, params_width));
   ram(166) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(80, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(725, params_width), to_signed(-1, params_width));
   ram(167) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(84, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(1052, params_width), to_signed(-1, params_width));
   ram(168) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(50, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(1225, params_width), to_signed(-1, params_width));
   ram(169) := ( to_signed(394, params_width), to_signed(2707802, params_width), to_signed(150, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(1262, params_width), to_signed(-1, params_width));
   ram(170) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(171) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(84, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(230, params_width), to_signed(0, params_width));
   ram(172) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(105, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(1195, params_width), to_signed(-1, params_width));
   ram(173) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(96, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-1678, params_width), to_signed(1, params_width));
   ram(174) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(59, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(-2219, params_width), to_signed(2, params_width));
   ram(175) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(112, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-3141, params_width), to_signed(2, params_width));
   ram(176) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(42, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-2007, params_width), to_signed(1, params_width));
   ram(177) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(64, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-4714, params_width), to_signed(3, params_width));
   ram(178) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(86, params_width), to_signed(-2, params_width), to_signed(-2, params_width), to_signed(4559, params_width), to_signed(-3, params_width));
   ram(179) := ( to_signed(390, params_width), to_signed(2835226, params_width), to_signed(110, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-3819, params_width), to_signed(3, params_width));
   ram(180) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(181) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(199, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(316, params_width), to_signed(0, params_width));
   ram(182) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(250, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-185, params_width), to_signed(0, params_width));
   ram(183) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(333, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(195, params_width), to_signed(0, params_width));
   ram(184) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(430, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(454, params_width), to_signed(0, params_width));
   ram(185) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(486, params_width), to_signed(2, params_width), to_signed(-2, params_width), to_signed(478, params_width), to_signed(-1, params_width));
   ram(186) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(615, params_width), to_signed(4, params_width), to_signed(-1, params_width), to_signed(-98, params_width), to_signed(0, params_width));
   ram(187) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(624, params_width), to_signed(18, params_width), to_signed(2, params_width), to_signed(1761, params_width), to_signed(-1, params_width));
   ram(188) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(850, params_width), to_signed(25, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(189) := ( to_signed(363, params_width), to_signed(2253, params_width), to_signed(1523, params_width), to_signed(32, params_width), to_signed(2, params_width), to_signed(2588, params_width), to_signed(-1, params_width));
   ram(190) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(191) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(192) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(107, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-354, params_width), to_signed(0, params_width));
   ram(193) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(85, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(1046, params_width), to_signed(-1, params_width));
   ram(194) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(120, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(5757, params_width), to_signed(-4, params_width));
   ram(195) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(120, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(8186, params_width), to_signed(-6, params_width));
   ram(196) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(73, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-2539, params_width), to_signed(2, params_width));
   ram(197) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(121, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-4685, params_width), to_signed(3, params_width));
   ram(198) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(114, params_width), to_signed(-2, params_width), to_signed(-2, params_width), to_signed(-1804, params_width), to_signed(1, params_width));
   ram(199) := ( to_signed(383, params_width), to_signed(2885171, params_width), to_signed(115, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-2236, params_width), to_signed(2, params_width));
   ram(200) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(201) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(124, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-727, params_width), to_signed(0, params_width));
   ram(202) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(133, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(200, params_width), to_signed(0, params_width));
   ram(203) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(114, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(321, params_width), to_signed(0, params_width));
   ram(204) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(112, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(980, params_width), to_signed(-1, params_width));
   ram(205) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(82, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(1138, params_width), to_signed(-1, params_width));
   ram(206) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(71, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(1441, params_width), to_signed(-1, params_width));
   ram(207) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(73, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(1858, params_width), to_signed(-1, params_width));
   ram(208) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(91, params_width), to_signed(-1, params_width), to_signed(-2, params_width), to_signed(1986, params_width), to_signed(-1, params_width));
   ram(209) := ( to_signed(361, params_width), to_signed(2961280, params_width), to_signed(142, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(2023, params_width), to_signed(-1, params_width));
   ram(210) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(211) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(212) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(219, params_width), to_signed(4, params_width), to_signed(0, params_width), to_signed(2263, params_width), to_signed(-1, params_width));
   ram(213) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(153, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(-5446, params_width), to_signed(3, params_width));
   ram(214) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(127, params_width), to_signed(-2, params_width), to_signed(-1, params_width), to_signed(-3197, params_width), to_signed(2, params_width));
   ram(215) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(79, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(-4703, params_width), to_signed(3, params_width));
   ram(216) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(24, params_width), to_signed(-3, params_width), to_signed(-2, params_width), to_signed(-624, params_width), to_signed(0, params_width));
   ram(217) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(-69, params_width), to_signed(-1, params_width), to_signed(-2, params_width), to_signed(493, params_width), to_signed(0, params_width));
   ram(218) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(-67, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(-18, params_width), to_signed(0, params_width));
   ram(219) := ( to_signed(433, params_width), to_signed(2898765, params_width), to_signed(-39, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(-4726, params_width), to_signed(3, params_width));
   ram(220) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(221) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(50, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(-376, params_width), to_signed(0, params_width));
   ram(222) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(85, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(1504, params_width), to_signed(-1, params_width));
   ram(223) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(80, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-7671, params_width), to_signed(5, params_width));
   ram(224) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(33, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(-947, params_width), to_signed(1, params_width));
   ram(225) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(114, params_width), to_signed(-6, params_width), to_signed(-1, params_width), to_signed(-1093, params_width), to_signed(1, params_width));
   ram(226) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(140, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(-1957, params_width), to_signed(1, params_width));
   ram(227) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(99, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(-432, params_width), to_signed(0, params_width));
   ram(228) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(93, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(2767, params_width), to_signed(-2, params_width));
   ram(229) := ( to_signed(193, params_width), to_signed(3202714, params_width), to_signed(327, params_width), to_signed(-3, params_width), to_signed(-3, params_width), to_signed(-5558, params_width), to_signed(3, params_width));
   ram(230) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(231) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(347, params_width), to_signed(0, params_width));
   ram(232) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(251, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(233) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-2655, params_width), to_signed(2, params_width));
   ram(234) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(235) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(162, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(236) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-5727, params_width), to_signed(3, params_width));
   ram(237) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(238) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(239) := ( to_signed(461, params_width), to_signed(3061, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(240) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(241) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(135, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-2472, params_width), to_signed(1, params_width));
   ram(242) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(133, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(-1679, params_width), to_signed(1, params_width));
   ram(243) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(135, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(-242, params_width), to_signed(0, params_width));
   ram(244) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(128, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-299, params_width), to_signed(0, params_width));
   ram(245) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(143, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-424, params_width), to_signed(0, params_width));
   ram(246) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(122, params_width), to_signed(1, params_width), to_signed(-2, params_width), to_signed(520, params_width), to_signed(0, params_width));
   ram(247) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(106, params_width), to_signed(-1, params_width), to_signed(-2, params_width), to_signed(1032, params_width), to_signed(-1, params_width));
   ram(248) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(112, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(686, params_width), to_signed(0, params_width));
   ram(249) := ( to_signed(358, params_width), to_signed(3167987, params_width), to_signed(176, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(478, params_width), to_signed(0, params_width));
   ram(250) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(251) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(275, params_width), to_signed(23, params_width), to_signed(-1, params_width), to_signed(145, params_width), to_signed(0, params_width));
   ram(252) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(354, params_width), to_signed(-4, params_width), to_signed(-1, params_width), to_signed(-394, params_width), to_signed(0, params_width));
   ram(253) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(438, params_width), to_signed(-3, params_width), to_signed(-1, params_width), to_signed(-703, params_width), to_signed(0, params_width));
   ram(254) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(460, params_width), to_signed(-14, params_width), to_signed(-2, params_width), to_signed(2110, params_width), to_signed(-1, params_width));
   ram(255) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(532, params_width), to_signed(5, params_width), to_signed(-2, params_width), to_signed(113, params_width), to_signed(0, params_width));
   ram(256) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(623, params_width), to_signed(-4, params_width), to_signed(-2, params_width), to_signed(-1595, params_width), to_signed(1, params_width));
   ram(257) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(810, params_width), to_signed(23, params_width), to_signed(0, params_width), to_signed(5680, params_width), to_signed(-4, params_width));
   ram(258) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(618, params_width), to_signed(27, params_width), to_signed(2, params_width), to_signed(949, params_width), to_signed(-1, params_width));
   ram(259) := ( to_signed(501, params_width), to_signed(2163, params_width), to_signed(529, params_width), to_signed(34, params_width), to_signed(5, params_width), to_signed(-38, params_width), to_signed(1, params_width));
   ram(260) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(261) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(141, params_width), to_signed(-3, params_width), to_signed(0, params_width), to_signed(-1707, params_width), to_signed(1, params_width));
   ram(262) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(121, params_width), to_signed(-7, params_width), to_signed(-1, params_width), to_signed(6787, params_width), to_signed(-4, params_width));
   ram(263) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(313, params_width), to_signed(-12, params_width), to_signed(-2, params_width), to_signed(-3650, params_width), to_signed(2, params_width));
   ram(264) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(306, params_width), to_signed(32, params_width), to_signed(0, params_width), to_signed(1800, params_width), to_signed(-1, params_width));
   ram(265) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(456, params_width), to_signed(-10, params_width), to_signed(-2, params_width), to_signed(-14022, params_width), to_signed(9, params_width));
   ram(266) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(188, params_width), to_signed(-32, params_width), to_signed(3, params_width), to_signed(6941, params_width), to_signed(-4, params_width));
   ram(267) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-23002, params_width), to_signed(14, params_width));
   ram(268) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(30668, params_width), to_signed(-19, params_width));
   ram(269) := ( to_signed(297, params_width), to_signed(2174, params_width), to_signed(1686, params_width), to_signed(50, params_width), to_signed(2, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(270) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(271) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(260, params_width), to_signed(0, params_width));
   ram(272) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(492, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-1918, params_width), to_signed(1, params_width));
   ram(273) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(465, params_width), to_signed(-5, params_width), to_signed(-1, params_width), to_signed(-2401, params_width), to_signed(1, params_width));
   ram(274) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(483, params_width), to_signed(-3, params_width), to_signed(-2, params_width), to_signed(-6534, params_width), to_signed(4, params_width));
   ram(275) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(473, params_width), to_signed(-5, params_width), to_signed(-2, params_width), to_signed(-5017, params_width), to_signed(3, params_width));
   ram(276) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(515, params_width), to_signed(8, params_width), to_signed(-2, params_width), to_signed(3814, params_width), to_signed(-2, params_width));
   ram(277) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(519, params_width), to_signed(10, params_width), to_signed(-1, params_width), to_signed(4846, params_width), to_signed(-3, params_width));
   ram(278) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(516, params_width), to_signed(11, params_width), to_signed(-1, params_width), to_signed(6020, params_width), to_signed(-3, params_width));
   ram(279) := ( to_signed(676, params_width), to_signed(1913, params_width), to_signed(889, params_width), to_signed(28, params_width), to_signed(2, params_width), to_signed(-6191, params_width), to_signed(4, params_width));
   ram(280) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(281) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(159, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-9, params_width), to_signed(0, params_width));
   ram(282) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(180, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-29, params_width), to_signed(0, params_width));
   ram(283) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(232, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-13, params_width), to_signed(0, params_width));
   ram(284) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(245, params_width), to_signed(3, params_width), to_signed(-1, params_width), to_signed(42, params_width), to_signed(0, params_width));
   ram(285) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(354, params_width), to_signed(1, params_width), to_signed(-1, params_width), to_signed(-103, params_width), to_signed(0, params_width));
   ram(286) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-779, params_width), to_signed(1, params_width));
   ram(287) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(-664, params_width), to_signed(1, params_width));
   ram(288) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(523, params_width), to_signed(-27, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(289) := ( to_signed(380, params_width), to_signed(3808, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(290) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(291) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(104, params_width), to_signed(1, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(0, params_width));
   ram(292) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(132, params_width), to_signed(3, params_width), to_signed(0, params_width), to_signed(-12, params_width), to_signed(0, params_width));
   ram(293) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(173, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-26, params_width), to_signed(0, params_width));
   ram(294) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(155, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(-13, params_width), to_signed(0, params_width));
   ram(295) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(167, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(12, params_width), to_signed(0, params_width));
   ram(296) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(170, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(52, params_width), to_signed(0, params_width));
   ram(297) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(260, params_width), to_signed(3, params_width), to_signed(-1, params_width), to_signed(-14, params_width), to_signed(0, params_width));
   ram(298) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(305, params_width), to_signed(6, params_width), to_signed(-1, params_width), to_signed(-83, params_width), to_signed(0, params_width));
   ram(299) := ( to_signed(341, params_width), to_signed(1704, params_width), to_signed(428, params_width), to_signed(8, params_width), to_signed(0, params_width), to_signed(142, params_width), to_signed(0, params_width));
   ram(300) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(0, params_width));
   ram(301) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(127, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(5, params_width), to_signed(0, params_width));
   ram(302) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(129, params_width), to_signed(0, params_width), to_signed(0, params_width), to_signed(25, params_width), to_signed(0, params_width));
   ram(303) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(124, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(35, params_width), to_signed(0, params_width));
   ram(304) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(133, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(61, params_width), to_signed(0, params_width));
   ram(305) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(141, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(56, params_width), to_signed(0, params_width));
   ram(306) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(139, params_width), to_signed(-1, params_width), to_signed(-1, params_width), to_signed(97, params_width), to_signed(0, params_width));
   ram(307) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(143, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(67, params_width), to_signed(0, params_width));
   ram(308) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(137, params_width), to_signed(0, params_width), to_signed(-2, params_width), to_signed(67, params_width), to_signed(0, params_width));
   ram(309) := ( to_signed(396, params_width), to_signed(2214810, params_width), to_signed(221, params_width), to_signed(0, params_width), to_signed(-1, params_width), to_signed(71, params_width), to_signed(0, params_width));
return ram;
end function;

end package body;