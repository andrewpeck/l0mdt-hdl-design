--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: rpc_z to 1st layer tube number 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library heg_roi_lib;
use heg_roi_lib.roi_types_pkg.all;

package roi_lut_BILA3 is

  -- add length of constant array
  constant ROM_BILA3_Z_MAX_SIZE : integer := 6550;

  constant ROI_BILA3_Z_MEM : roi_z_lut_t(0 to ROM_BILA3_Z_MAX_SIZE - 1) := (

    0 to 329 => -1,
    330 to 359 =>0,
    360 to 389 =>1,
    390 to 419 =>2,
    420 to 449 =>3,
    450 to 479 =>4,
    480 to 509 =>5,
    510 to 539 =>6,
    540 to 569 =>7,
    570 to 599 =>8,
    600 to 629 =>9,
    630 to 659 =>10,
    660 to 689 =>11,
    690 to 719 =>12,
    720 to 749 =>13,
    750 to 779 =>14,
    780 to 809 =>15,
    810 to 838 =>16,
    839 to 868 =>17,
    869 to 898 =>18,
    899 to 928 =>19,
    929 to 958 =>20,
    959 to 988 =>21,
    989 to 1018 =>22,
    1019 to 1048 =>23,
    1049 to 1078 =>24,
    1079 to 1108 =>25,
    1109 to 1138 =>26,
    1139 to 1168 =>27,
    1169 to 1198 =>28,
    1199 to 1228 =>29,
    1229 to 1249 =>-1,
    1250 to 1279 =>30,
    1280 to 1309 =>31,
    1310 to 1339 =>32,
    1340 to 1369 =>33,
    1370 to 1399 =>34,
    1400 to 1429 =>35,
    1430 to 1459 =>36,
    1460 to 1489 =>37,
    1490 to 1519 =>38,
    1520 to 1549 =>39,
    1550 to 1579 =>40,
    1580 to 1609 =>41,
    1610 to 1639 =>42,
    1640 to 1669 =>43,
    1670 to 1699 =>44,
    1700 to 1729 =>45,
    1730 to 1758 =>46,
    1759 to 1788 =>47,
    1789 to 1818 =>48,
    1819 to 1848 =>49,
    1849 to 1878 =>50,
    1879 to 1908 =>51,
    1909 to 1938 =>52,
    1939 to 1968 =>53,
    1969 to 1998 =>54,
    1999 to 2028 =>55,
    2029 to 2058 =>56,
    2059 to 2088 =>57,
    2089 to 2118 =>58,
    2119 to 2148 =>59,
    2149 to 2178 =>60,
    2179 to 2208 =>61,
    2209 to 2238 =>62,
    2239 to 2268 =>63,
    2269 to 2298 =>64,
    2299 to 2328 =>65,
    2329 to 2349 =>-1,
    2350 to 2379 =>66,
    2380 to 2409 =>67,
    2410 to 2439 =>68,
    2440 to 2469 =>69,
    2470 to 2499 =>70,
    2500 to 2529 =>71,
    2530 to 2559 =>72,
    2560 to 2589 =>73,
    2590 to 2619 =>74,
    2620 to 2649 =>75,
    2650 to 2679 =>76,
    2680 to 2709 =>77,
    2710 to 2739 =>78,
    2740 to 2769 =>79,
    2770 to 2799 =>80,
    2800 to 2829 =>81,
    2830 to 2858 =>82,
    2859 to 2888 =>83,
    2889 to 2918 =>84,
    2919 to 2948 =>85,
    2949 to 2978 =>86,
    2979 to 3008 =>87,
    3009 to 3038 =>88,
    3039 to 3068 =>89,
    3069 to 3098 =>90,
    3099 to 3128 =>91,
    3129 to 3158 =>92,
    3159 to 3188 =>93,
    3189 to 3218 =>94,
    3219 to 3248 =>95,
    3249 to 3449 =>-1,
    3450 to 3479 =>96,
    3480 to 3509 =>97,
    3510 to 3539 =>98,
    3540 to 3569 =>99,
    3570 to 3599 =>100,
    3600 to 3629 =>101,
    3630 to 3659 =>102,
    3660 to 3689 =>103,
    3690 to 3719 =>104,
    3720 to 3749 =>105,
    3750 to 3779 =>106,
    3780 to 3809 =>107,
    3810 to 3839 =>108,
    3840 to 3869 =>109,
    3870 to 3899 =>110,
    3900 to 3929 =>111,
    3930 to 3958 =>112,
    3959 to 3988 =>113,
    3989 to 4018 =>114,
    4019 to 4048 =>115,
    4049 to 4078 =>116,
    4079 to 4108 =>117,
    4109 to 4138 =>118,
    4139 to 4168 =>119,
    4169 to 4198 =>120,
    4199 to 4228 =>121,
    4229 to 4258 =>122,
    4259 to 4288 =>123,
    4289 to 4318 =>124,
    4319 to 4348 =>125,
    4349 to 4378 =>126,
    4379 to 4408 =>127,
    4409 to 4438 =>128,
    4439 to 4468 =>129,
    4469 to 4498 =>130,
    4499 to 4528 =>131,
    4529 to 4549 =>-1,
    4550 to 4579 =>132,
    4580 to 4609 =>133,
    4610 to 4639 =>134,
    4640 to 4669 =>135,
    4670 to 4699 =>136,
    4700 to 4729 =>137,
    4730 to 4759 =>138,
    4760 to 4789 =>139,
    4790 to 4819 =>140,
    4820 to 4849 =>141,
    4850 to 4879 =>142,
    4880 to 4909 =>143,
    4910 to 4939 =>144,
    4940 to 4969 =>145,
    4970 to 4999 =>146,
    5000 to 5029 =>147,
    5030 to 5058 =>148,
    5059 to 5088 =>149,
    5089 to 5118 =>150,
    5119 to 5148 =>151,
    5149 to 5178 =>152,
    5179 to 5208 =>153,
    5209 to 5238 =>154,
    5239 to 5268 =>155,
    5269 to 5298 =>156,
    5299 to 5328 =>157,
    5329 to 5358 =>158,
    5359 to 5388 =>159,
    5389 to 5418 =>160,
    5419 to 5448 =>161,
    5449 to 5469 =>-1,
    5470 to 5499 =>162,
    5500 to 5529 =>163,
    5530 to 5559 =>164,
    5560 to 5589 =>165,
    5590 to 5619 =>166,
    5620 to 5649 =>167,
    5650 to 5679 =>168,
    5680 to 5709 =>169,
    5710 to 5739 =>170,
    5740 to 5769 =>171,
    5770 to 5799 =>172,
    5800 to 5829 =>173,
    5830 to 5859 =>174,
    5860 to 5889 =>175,
    5890 to 5919 =>176,
    5920 to 5949 =>177,
    5950 to 5978 =>178,
    5979 to 6008 =>179,
    6009 to 6038 =>180,
    6039 to 6068 =>181,
    6069 to 6098 =>182,
    6099 to 6128 =>183,
    6129 to 6158 =>184,
    6159 to 6188 =>185,
    6189 to 6218 =>186,
    6219 to 6248 =>187,
    6249 to 6278 =>188,
    6279 to 6308 =>189,
    6309 to 6338 =>190,
    6339 to 6368 =>191,
    6369 to 6398 =>192,
    6399 to 6428 =>193,
    6429 to 6458 =>194,
    6459 to 6488 =>195,
    6489 to 6518 =>196,
    6519 to 6549 =>197
  );

 end package roi_lut_BILA3;
