--------------------------------------------------------------------------------
-- UMass , Physics Department
-- Project: ult
-- File: top_ult_sim.vhd
-- Module: <<moduleName>>
-- File PATH: /top_ult_sim.vhd
-- -----
-- File Created: Wednesday, 8th June 2022 9:54:45 am
-- Author: Guillermo Loustau de Linares (guillermo.ldl@cern.ch)
-- -----
-- Last Modified: Saturday, 11th February 2023 12:49:28 am
-- Modified By: Guillermo Loustau de Linares (guillermo.ldl@cern.ch>)
-- -----
-- HISTORY:
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_misc.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;
use shared_lib.config_pkg.all;
-- use shared_lib.vhdl2008_functions_pkg.all;
use shared_lib.detector_param_pkg.all;

library ult_lib;

library ctrl_lib;
use ctrl_lib.HPS_CTRL.all;
use ctrl_lib.TAR_CTRL.all;
use ctrl_lib.MTC_CTRL.all;
use ctrl_lib.UCM_CTRL.all;
use ctrl_lib.DAQ_CTRL.all;
use ctrl_lib.TF_CTRL.all;
use ctrl_lib.MPL_CTRL.all;
use ctrl_lib.FM_CTRL.all;

library fm_lib;
use fm_lib.fm_ult_pkg.all;

entity ult_tb is
  port (
    PRJ_INFO            : string  := "not_defined";
    IN_SLC_FILE         : string  := "not_defined.csv";
    IN_CTRL_FILE        : string  := "not_defined.csv";
    DUMMY               : boolean := false
  );
end entity ult_tb;

architecture beh of ult_tb is
  signal clock_and_control     : l0mdt_control_rt;

  signal i_inner_tdc_hits  : tdcpolmux2tar_avt (c_HPS_MAX_HP_INN -1 downto 0);
  signal i_middle_tdc_hits : tdcpolmux2tar_avt (c_HPS_MAX_HP_MID -1 downto 0);
  signal i_outer_tdc_hits  : tdcpolmux2tar_avt (c_HPS_MAX_HP_OUT -1 downto 0);
  signal i_extra_tdc_hits  : tdcpolmux2tar_avt (c_HPS_MAX_HP_EXT -1 downto 0);

  signal i_main_primary_slc        :slc_rx_avt(2 downto 0);  -- is the main SL used
  signal i_main_secondary_slc      :slc_rx_avt(2 downto 0);  -- only used in the big endcap
  signal i_plus_neighbor_slc       :slc_rx_vt;
  signal i_minus_neighbor_slc      :slc_rx_vt;

  signal i_plus_neighbor_segments  : sf2ptcalc_avt(c_NUM_SF_INPUTS - 1 downto 0);
  signal i_minus_neighbor_segments : sf2ptcalc_avt(c_NUM_SF_INPUTS - 1 downto 0);

  signal hps_inn_ctrl_r        : HPS_CTRL_t;
  signal hps_inn_mon_r         : HPS_MON_t;
  signal hps_mid_ctrl_r        : HPS_CTRL_t;
  signal hps_mid_mon_r         : HPS_MON_t;
  signal hps_out_ctrl_r        : HPS_CTRL_t;
  signal hps_out_mon_r         : HPS_MON_t;
  signal hps_ext_ctrl_r        : HPS_CTRL_t;
  signal hps_ext_mon_r         : HPS_MON_t;

  signal tar_inn_ctrl_r        : TAR_CTRL_t;
  signal tar_inn_mon_r         : TAR_MON_t;
  signal tar_mid_ctrl_r        : TAR_CTRL_t;
  signal tar_mid_mon_r         : TAR_MON_t;
  signal tar_out_ctrl_r        : TAR_CTRL_t;
  signal tar_out_mon_r         : TAR_MON_t;
  signal tar_ext_ctrl_r        : TAR_CTRL_t;
  signal tar_ext_mon_r         : TAR_MON_t;

  signal mtc_ctrl_r            : MTC_CTRL_t;
  signal mtc_mon_r             : MTC_MON_t;
  signal ucm_ctrl_r            : UCM_CTRL_t;
  signal ucm_mon_r             : UCM_MON_t;
  signal daq_ctrl_r            : DAQ_CTRL_t;
  signal daq_mon_r             : DAQ_MON_t;
  signal tf_ctrl_r             : TF_CTRL_t;
  signal tf_mon_r              : TF_MON_t;
  signal mpl_ctrl_r            : MPL_CTRL_t;
  signal mpl_mon_r             : MPL_MON_t;
  signal fm_ctrl_r             : FM_CTRL_t;
  signal fm_mon_r              : FM_MON_t;

  signal hps_inn_ctrl_v        : std_logic_vector(HPS_CTRL_t'w -1 downto 0); -- : in  H2S_CTRL_t;
  signal hps_inn_mon_v         : std_logic_vector(HPS_MON_t'w -1 downto 0);--  : out H2S_MON_t;
  signal hps_mid_ctrl_v        : std_logic_vector(HPS_CTRL_t'w -1 downto 0); -- : in  H2S_CTRL_t;
  signal hps_mid_mon_v         : std_logic_vector(HPS_MON_t'w -1 downto 0);--  : out H2S_MON_t;
  signal hps_out_ctrl_v        : std_logic_vector(HPS_CTRL_t'w -1 downto 0); -- : in  H2S_CTRL_t;
  signal hps_out_mon_v         : std_logic_vector(HPS_MON_t'w -1 downto 0);--  : out H2S_MON_t;
  signal hps_ext_ctrl_v        : std_logic_vector(HPS_CTRL_t'w -1 downto 0); -- : in  H2S_CTRL_t;
  signal hps_ext_mon_v         : std_logic_vector(HPS_MON_t'w -1 downto 0);--  : out H2S_MON_t;
  
  signal tar_inn_ctrl_v        : std_logic_vector(TAR_CTRL_t'w -1 downto 0);
  signal tar_inn_mon_v         : std_logic_vector(TAR_MON_t'w -1 downto 0);
  signal tar_mid_ctrl_v        : std_logic_vector(TAR_CTRL_t'w -1 downto 0);
  signal tar_mid_mon_v         : std_logic_vector(TAR_MON_t'w -1 downto 0);
  signal tar_out_ctrl_v        : std_logic_vector(TAR_CTRL_t'w -1 downto 0);
  signal tar_out_mon_v         : std_logic_vector(TAR_MON_t'w -1 downto 0);
  signal tar_ext_ctrl_v        : std_logic_vector(TAR_CTRL_t'w -1 downto 0);
  signal tar_ext_mon_v         : std_logic_vector(TAR_MON_t'w -1 downto 0);

  signal mtc_ctrl_v            : std_logic_vector(MTC_CTRL_t'w -1 downto 0);
  signal mtc_mon_v             : std_logic_vector(MTC_MON_t'w -1 downto 0);

  signal ucm_ctrl_v            : std_logic_vector(UCM_CTRL_t'w -1 downto 0);
  signal ucm_mon_v             : std_logic_vector(UCM_MON_t'w -1 downto 0);
  
  signal daq_ctrl_v            : std_logic_vector(DAQ_CTRL_t'w -1 downto 0);
  signal daq_mon_v             : std_logic_vector(DAQ_MON_t'w -1 downto 0);
  
  signal tf_ctrl_v             : std_logic_vector(TF_CTRL_t'w -1 downto 0);
  signal tf_mon_v              : std_logic_vector(TF_MON_t'w -1 downto 0);
  
  signal mpl_ctrl_v            : std_logic_vector(MPL_CTRL_t'w -1 downto 0);
  signal mpl_mon_v             : std_logic_vector(MPL_MON_t'w -1 downto 0);
  
  signal fm_ctrl_v             : std_logic_vector(FM_CTRL_t'w -1 downto 0);
  signal fm_mon_v              : std_logic_vector(FM_MON_t'w -1 downto 0);

  signal o_daq_streams     : felix_stream_avt (c_DAQ_LINKS - 1 downto 0);

  signal o_plus_neighbor_segments  : sf2ptcalc_avt(c_NUM_SF_OUTPUTS - 1 downto 0);
  signal o_minus_neighbor_segments : sf2ptcalc_avt(c_NUM_SF_OUTPUTS - 1 downto 0);

  signal o_MTC : mtc_out_avt(c_NUM_MTC-1 downto 0);
  signal o_NSP : mtc2nsp_avt(c_NUM_NSP-1 downto 0);

begin
  
  ULT : entity ult_lib.ult
  generic map(
    DUMMY       => DUMMY
    )
  port map(
    -- pipeline clock
    clock_and_control => clock_and_control,
    ttc_commands      => ttc_commands,

    -- TDC Hits from Polmux
    i_inn_tdc_hits_av => i_inner_tdc_hits,
    i_mid_tdc_hits_av => i_middle_tdc_hits,
    i_out_tdc_hits_av => i_outer_tdc_hits,
    i_ext_tdc_hits_av => i_extra_tdc_hits,

    -- TAR Hits for simulation
    -- i_inner_tar_hits  => i_inner_tar_hits,
    -- i_middle_tar_hits => i_middle_tar_hits,
    -- i_outer_tar_hits  => i_outer_tar_hits,
    -- i_extra_tar_hits  => i_extra_tar_hits,

    -- Sector Logic Candidates
    i_main_primary_slc   => i_main_primary_slc,
    i_main_secondary_slc => i_main_secondary_slc,
    i_plus_neighbor_slc  => i_plus_neighbor_slc,
    i_minus_neighbor_slc => i_minus_neighbor_slc,

    -- Segments in from neighbor
    i_plus_neighbor_segments  => i_plus_neighbor_segments,
    i_minus_neighbor_segments => i_minus_neighbor_segments,

    -- ULT Control

    hps_inn_ctrl_v => hps_inn_ctrl_v ,
    hps_inn_mon_v  => hps_inn_mon_v  ,
    hps_mid_ctrl_v => hps_mid_ctrl_v ,
    hps_mid_mon_v  => hps_mid_mon_v  ,
    hps_out_ctrl_v => hps_out_ctrl_v ,
    hps_out_mon_v  => hps_out_mon_v  ,
    hps_ext_ctrl_v => hps_ext_ctrl_v ,
    hps_ext_mon_v  => hps_ext_mon_v  ,
    tar_inn_ctrl_v => tar_inn_ctrl_v,
    tar_inn_mon_v  => tar_inn_mon_v ,
    tar_mid_ctrl_v => tar_mid_ctrl_v,
    tar_mid_mon_v  => tar_mid_mon_v ,
    tar_out_ctrl_v => tar_out_ctrl_v,
    tar_out_mon_v  => tar_out_mon_v ,
    tar_ext_ctrl_v => tar_ext_ctrl_v,
    tar_ext_mon_v  => tar_ext_mon_v ,
    mtc_ctrl_v => mtc_ctrl_v,
    mtc_mon_v  => mtc_mon_v,
    ucm_ctrl_v => ucm_ctrl_v,
    ucm_mon_v  => ucm_mon_v,
    daq_ctrl_v => daq_ctrl_v,
    daq_mon_v  => daq_mon_v,
    tf_ctrl_v  => tf_ctrl_v,
    tf_mon_v   => tf_mon_v,
    mpl_ctrl_v => mpl_ctrl_v,
    mpl_mon_v  => mpl_mon_v,
    fm_ctrl_v  => fm_ctrl_v,
    fm_mon_v   => fm_mon_v,

    
    -- Array of DAQ data streams (e.g. 64 bit strams) to send to MGT
    o_daq_streams => o_daq_streams,

    -- Segments Out to Neighbor
    o_plus_neighbor_segments_av  => o_plus_neighbor_segments,
    o_minus_neighbor_segments_av => o_minus_neighbor_segments,

    -- MUCTPI
    o_MTC => o_MTC,
    o_NSP => o_NSP,

    sump => sump
);
  
  
end architecture beh;



-- entity top_ult is
--   generic (
--     DUMMY       : boolean := false

--     -- g_h2s_ctrl  : H2S_CTRL_t := zero(g_h2s_ctrl);
--     );

--   port (
--     -- pipeline clock
--     -- clock_and_control : in l0mdt_control_rt;
--     clk                 : in std_logic;
--     rst                 : in std_logic;
--     bx                  : in std_logic;

--     ttc_commands        : in l0mdt_ttc_rt;

--     -- axi control

--     h2s_ctrl_r            : in  H2S_CTRL_t;
--     h2s_mon_r             : out H2S_MON_t;

--     tar_ctrl_r            : in  TAR_CTRL_t;
--     tar_mon_r             : out TAR_MON_t;

--     mtc_ctrl_r            : in  MTC_CTRL_t;
--     mtc_mon_r             : out MTC_MON_t;

--     ucm_ctrl_r            : in  UCM_CTRL_t;
--     ucm_mon_r             : out UCM_MON_t;

--     daq_ctrl_r            : in  DAQ_CTRL_t;
--     daq_mon_r             : out DAQ_MON_t;

--     tf_ctrl_r             : in  TF_CTRL_t;
--     tf_mon_r              : out TF_MON_t;

--     mpl_ctrl_r            : in  MPL_CTRL_t;
--     mpl_mon_r             : out MPL_MON_t;

--     fm_ctrl_r             : in FM_CTRL_t;
--     fm_mon_r              : out FM_MON_t;

--     -- TDC Hits from Polmux
--     i_inner_tdc_hits  : in tdcpolmux2tar_avt (c_HPS_MAX_HP_INN -1 downto 0);
--     i_middle_tdc_hits : in tdcpolmux2tar_avt (c_HPS_MAX_HP_MID -1 downto 0);
--     i_outer_tdc_hits  : in tdcpolmux2tar_avt (c_HPS_MAX_HP_OUT -1 downto 0);
--     i_extra_tdc_hits  : in tdcpolmux2tar_avt (c_HPS_MAX_HP_EXT -1 downto 0);

--     -- TDC Hits from Tar
--     -- i_inner_tar_hits  : in tar2hps_avt (c_EN_TAR_HITS*c_HPS_MAX_HP_INN -1 downto 0);
--     -- i_middle_tar_hits : in tar2hps_avt (c_EN_TAR_HITS*c_HPS_MAX_HP_MID -1 downto 0);
--     -- i_outer_tar_hits  : in tar2hps_avt (c_EN_TAR_HITS*c_HPS_MAX_HP_OUT -1 downto 0);
--     -- i_extra_tar_hits  : in tar2hps_avt (c_EN_TAR_HITS*c_HPS_MAX_HP_EXT -1 downto 0);

--     -- Sector Logic Candidates
--     i_main_primary_slc        : in slc_rx_avt(2 downto 0);  -- is the main SL used
--     i_main_secondary_slc      : in slc_rx_avt(2 downto 0);  -- only used in the big endcap
--     i_plus_neighbor_slc       : in slc_rx_vt;
--     i_minus_neighbor_slc      : in slc_rx_vt;
--     -- Segments in from neighbor
--     i_plus_neighbor_segments  : in sf2ptcalc_avt(c_NUM_SF_INPUTS - 1 downto 0);
--     i_minus_neighbor_segments : in sf2ptcalc_avt(c_NUM_SF_INPUTS - 1 downto 0);

--     -- Array of DAQ data streams (e.g. 64 bit strams) to send to MGT
--     o_daq_streams     : out felix_stream_avt (c_HPS_MAX_HP_INN
--                                                   + c_HPS_MAX_HP_MID
--                                                   + c_HPS_MAX_HP_OUT - 1 downto 0);
--     -- o_daq_streams : out felix_stream_avt (c_NUM_DAQ_STREAMS-1 downto 0);

--     -- Segments Out to Neighbor
--     o_plus_neighbor_segments  : out sf2ptcalc_avt(c_NUM_SF_OUTPUTS - 1 downto 0);
--     o_minus_neighbor_segments : out sf2ptcalc_avt(c_NUM_SF_OUTPUTS - 1 downto 0);

--     -- MUCTPI
--     o_MTC : out mtc_out_avt(c_NUM_MTC-1 downto 0);
--     o_NSP : out mtc2nsp_avt(c_NUM_NSP-1 downto 0);

--     sump : out std_logic

--     );

-- end entity top_ult;

-- architecture behavioral of top_ult is
--   signal clock_and_control : l0mdt_control_rt;

--   signal h2s_ctrl_v            : std_logic_vector(len(h2s_ctrl_r ) -1 downto 0);
--   signal h2s_mon_v             : std_logic_vector(len(h2s_mon_r  ) -1 downto 0);
--   signal tar_ctrl_v            : std_logic_vector(len(tar_ctrl_r ) -1 downto 0);
--   signal tar_mon_v             : std_logic_vector(len(tar_mon_r  ) -1 downto 0);
--   signal mtc_ctrl_v            : std_logic_vector(len(mtc_ctrl_r ) -1 downto 0);
--   signal mtc_mon_v             : std_logic_vector(len(mtc_mon_r  ) -1 downto 0);
--   signal ucm_ctrl_v            : std_logic_vector(len(ucm_ctrl_r ) -1 downto 0);
--   signal ucm_mon_v             : std_logic_vector(len(ucm_mon_r  ) -1 downto 0);
--   signal daq_ctrl_v            : std_logic_vector(len(daq_ctrl_r ) -1 downto 0);
--   signal daq_mon_v             : std_logic_vector(len(daq_mon_r  ) -1 downto 0);
--   signal tf_ctrl_v             : std_logic_vector(len(tf_ctrl_r  ) -1 downto 0);
--   signal tf_mon_v              : std_logic_vector(len(tf_mon_r   ) -1 downto 0);
--   signal mpl_ctrl_v            : std_logic_vector(len(mpl_ctrl_r ) -1 downto 0);
--   signal mpl_mon_v             : std_logic_vector(len(mpl_mon_r  ) -1 downto 0);
--   signal fm_ctrl_v             : std_logic_vector(len(fm_ctrl_r  ) -1 downto 0);
--   signal fm_mon_v              : std_logic_vector(len(fm_mon_r  ) -1 downto 0);
-- begin

--   -- ctrl/mon
--   ucm_ctrl_v  <= convert(ucm_ctrl_r,ucm_ctrl_v);
--   ucm_mon_r   <= convert(ucm_mon_v,ucm_mon_r);
--   tar_ctrl_v  <= convert(tar_ctrl_r,tar_ctrl_v);
--   tar_mon_r   <= convert(tar_mon_v,tar_mon_r);
--   h2s_ctrl_v  <= convert(h2s_ctrl_r,h2s_ctrl_v);
--   h2s_mon_r   <= convert(h2s_mon_v,h2s_mon_r);
--   mpl_ctrl_v  <= convert(mpl_ctrl_r,mpl_ctrl_v);
--   mpl_mon_r   <= convert(mpl_mon_v,mpl_mon_r);
--   tf_ctrl_v   <= convert(tf_ctrl_r,tf_ctrl_v);
--   tf_mon_r    <= convert(tf_mon_v,tf_mon_r);
--   mtc_ctrl_v  <= convert(mtc_ctrl_r,mtc_ctrl_v);
--   mtc_mon_r   <= convert(mtc_mon_v,mtc_mon_r);
--   daq_ctrl_v  <= convert(daq_ctrl_r,daq_ctrl_v);
--   daq_mon_r   <= convert(daq_mon_v,daq_mon_r);
--   fm_ctrl_v   <= convert(fm_ctrl_r,fm_ctrl_v);
--   fm_mon_r    <= convert(fm_mon_v,fm_mon_r);
  
  
--   clock_and_control.clk <= clk;
--   clock_and_control.rst <= rst;
--   clock_and_control.bx  <= bx;


--   ULT : entity ult_lib.ult
--     generic map(
--       DUMMY       => DUMMY
--       )
--     port map(
--       -- pipeline clock
--       clock_and_control => clock_and_control,
--       ttc_commands      => ttc_commands,

--       -- TDC Hits from Polmux
--       i_inn_tdc_hits_av => i_inner_tdc_hits,
--       i_mid_tdc_hits_av => i_middle_tdc_hits,
--       i_out_tdc_hits_av => i_outer_tdc_hits,
--       i_ext_tdc_hits_av => i_extra_tdc_hits,

--       -- TAR Hits for simulation
--       -- i_inner_tar_hits  => i_inner_tar_hits,
--       -- i_middle_tar_hits => i_middle_tar_hits,
--       -- i_outer_tar_hits  => i_outer_tar_hits,
--       -- i_extra_tar_hits  => i_extra_tar_hits,

--       -- Sector Logic Candidates
--       i_main_primary_slc   => i_main_primary_slc,
--       i_main_secondary_slc => i_main_secondary_slc,
--       i_plus_neighbor_slc  => i_plus_neighbor_slc,
--       i_minus_neighbor_slc => i_minus_neighbor_slc,

--       -- Segments in from neighbor
--       i_plus_neighbor_segments  => i_plus_neighbor_segments,
--       i_minus_neighbor_segments => i_minus_neighbor_segments,

--       -- ULT Control

--       h2s_ctrl_v => h2s_ctrl_v,
--       h2s_mon_v  => h2s_mon_v,
--       tar_ctrl_v => tar_ctrl_v,
--       tar_mon_v  => tar_mon_v,
--       mtc_ctrl_v => mtc_ctrl_v,
--       mtc_mon_v  => mtc_mon_v,
--       ucm_ctrl_v => ucm_ctrl_v,
--       ucm_mon_v  => ucm_mon_v,
--       daq_ctrl_v => daq_ctrl_v,
--       daq_mon_v  => daq_mon_v,
--       tf_ctrl_v  => tf_ctrl_v,
--       tf_mon_v   => tf_mon_v,
--       mpl_ctrl_v => mpl_ctrl_v,
--       mpl_mon_v  => mpl_mon_v,

--       fm_ctrl_v  => fm_ctrl_v,
--       fm_mon_v   => fm_mon_v,

--       -- Array of DAQ data streams (e.g. 64 bit strams) to send to MGT
--       o_daq_streams => o_daq_streams,

--       -- Segments Out to Neighbor
--       o_plus_neighbor_segments_av  => o_plus_neighbor_segments,
--       o_minus_neighbor_segments_av => o_minus_neighbor_segments,

--       -- MUCTPI
--       o_MTC => o_MTC,
--       o_NSP => o_NSP,

--       sump => sump
--       );


-- end behavioral;
