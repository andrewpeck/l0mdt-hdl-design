library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library shared_lib;
use shared_lib.interfaces_types.all;

package ucm_pkg is

end package ucm_pkg;


------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package body ucm_pkg is

end package body ucm_pkg;
