--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: angle (mrad) to slope 
--  Slope multiplier: 1024 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package roi_tan is

    -- add length of constant array
    constant ROM_TAN_MAX_SIZE : integer := 1569;
    type roi_tan_lut_t is array (integer range <>) of integer;

    constant ROI_TAN_MEM : roi_tan_lut_t(0 to ROM_TAN_MAX_SIZE - 1) := (

       0  => 1024003,
       1  => 512000,
       2  => 341333,
       3  => 255999,
       4  => 204798,
       5  => 170665,
       6  => 146283,
       7  => 127997,
       8  => 113775,
       9  => 102397,
      10  => 93087,
      11  => 85329,
      12  => 78765,
      13  => 73138,
      14  => 68262,
      15  => 63995,
      16  => 60230,
      17  => 56883,
      18  => 53888,
      19  => 51193,
      20  => 48755,
      21  => 46538,
      22  => 44514,
      23  => 42658,
      24  => 40951,
      25  => 39376,
      26  => 37917,
      27  => 36562,
      28  => 35300,
      29  => 34123,
      30  => 33022,
      31  => 31989,
      32  => 31019,
      33  => 30106,
      34  => 29245,
      35  => 28432,
      36  => 27663,
      37  => 26934,
      38  => 26243,
      39  => 25586,
      40  => 24962,
      41  => 24367,
      42  => 23799,
      43  => 23258,
      44  => 22740,
      45  => 22245,
      46  => 21771,
      47  => 21317,
      48  => 20881,
      49  => 20463,
      50  => 20061,
      51  => 19675,
      52  => 19303,
      53  => 18945,
      54  => 18599,
      55  => 18267,
      56  => 17945,
      57  => 17635,
      58  => 17336,
      59  => 17046,
      60  => 16766,
      61  => 16495,
      62  => 16232,
      63  => 15978,
      64  => 15732,
      65  => 15493,
      66  => 15261,
      67  => 15036,
      68  => 14817,
      69  => 14605,
      70  => 14398,
      71  => 14198,
      72  => 14002,
      73  => 13813,
      74  => 13628,
      75  => 13448,
      76  => 13272,
      77  => 13102,
      78  => 12935,
      79  => 12773,
      80  => 12614,
      81  => 12460,
      82  => 12309,
      83  => 12162,
      84  => 12018,
      85  => 11878,
      86  => 11740,
      87  => 11606,
      88  => 11475,
      89  => 11347,
      90  => 11222,
      91  => 11099,
      92  => 10979,
      93  => 10862,
      94  => 10747,
      95  => 10634,
      96  => 10524,
      97  => 10416,
      98  => 10310,
      99  => 10206,
     100  => 10104,
     101  => 10004,
     102  =>  9907,
     103  =>  9811,
     104  =>  9717,
     105  =>  9624,
     106  =>  9534,
     107  =>  9445,
     108  =>  9357,
     109  =>  9272,
     110  =>  9187,
     111  =>  9105,
     112  =>  9023,
     113  =>  8944,
     114  =>  8865,
     115  =>  8788,
     116  =>  8712,
     117  =>  8638,
     118  =>  8564,
     119  =>  8492,
     120  =>  8421,
     121  =>  8352,
     122  =>  8283,
     123  =>  8216,
     124  =>  8149,
     125  =>  8084,
     126  =>  8020,
     127  =>  7956,
     128  =>  7894,
     129  =>  7832,
     130  =>  7772,
     131  =>  7712,
     132  =>  7654,
     133  =>  7596,
     134  =>  7539,
     135  =>  7483,
     136  =>  7428,
     137  =>  7373,
     138  =>  7319,
     139  =>  7266,
     140  =>  7214,
     141  =>  7163,
     142  =>  7112,
     143  =>  7062,
     144  =>  7013,
     145  =>  6964,
     146  =>  6916,
     147  =>  6868,
     148  =>  6822,
     149  =>  6775,
     150  =>  6730,
     151  =>  6685,
     152  =>  6641,
     153  =>  6597,
     154  =>  6553,
     155  =>  6511,
     156  =>  6469,
     157  =>  6427,
     158  =>  6386,
     159  =>  6345,
     160  =>  6305,
     161  =>  6266,
     162  =>  6226,
     163  =>  6188,
     164  =>  6150,
     165  =>  6112,
     166  =>  6075,
     167  =>  6038,
     168  =>  6001,
     169  =>  5965,
     170  =>  5930,
     171  =>  5895,
     172  =>  5860,
     173  =>  5826,
     174  =>  5792,
     175  =>  5758,
     176  =>  5725,
     177  =>  5692,
     178  =>  5659,
     179  =>  5627,
     180  =>  5596,
     181  =>  5564,
     182  =>  5533,
     183  =>  5502,
     184  =>  5472,
     185  =>  5442,
     186  =>  5412,
     187  =>  5382,
     188  =>  5353,
     189  =>  5324,
     190  =>  5296,
     191  =>  5268,
     192  =>  5240,
     193  =>  5212,
     194  =>  5185,
     195  =>  5157,
     196  =>  5131,
     197  =>  5104,
     198  =>  5078,
     199  =>  5052,
     200  =>  5026,
     201  =>  5000,
     202  =>  4975,
     203  =>  4950,
     204  =>  4925,
     205  =>  4900,
     206  =>  4876,
     207  =>  4852,
     208  =>  4828,
     209  =>  4804,
     210  =>  4781,
     211  =>  4758,
     212  =>  4735,
     213  =>  4712,
     214  =>  4689,
     215  =>  4667,
     216  =>  4645,
     217  =>  4623,
     218  =>  4601,
     219  =>  4579,
     220  =>  4558,
     221  =>  4537,
     222  =>  4516,
     223  =>  4495,
     224  =>  4474,
     225  =>  4454,
     226  =>  4433,
     227  =>  4413,
     228  =>  4393,
     229  =>  4373,
     230  =>  4354,
     231  =>  4334,
     232  =>  4315,
     233  =>  4296,
     234  =>  4277,
     235  =>  4258,
     236  =>  4239,
     237  =>  4221,
     238  =>  4203,
     239  =>  4184,
     240  =>  4166,
     241  =>  4148,
     242  =>  4131,
     243  =>  4113,
     244  =>  4096,
     245  =>  4078,
     246  =>  4061,
     247  =>  4044,
     248  =>  4027,
     249  =>  4010,
     250  =>  3994,
     251  =>  3977,
     252  =>  3961,
     253  =>  3944,
     254  =>  3928,
     255  =>  3912,
     256  =>  3896,
     257  =>  3881,
     258  =>  3865,
     259  =>  3849,
     260  =>  3834,
     261  =>  3819,
     262  =>  3803,
     263  =>  3788,
     264  =>  3773,
     265  =>  3758,
     266  =>  3744,
     267  =>  3729,
     268  =>  3714,
     269  =>  3700,
     270  =>  3686,
     271  =>  3671,
     272  =>  3657,
     273  =>  3643,
     274  =>  3629,
     275  =>  3615,
     276  =>  3602,
     277  =>  3588,
     278  =>  3575,
     279  =>  3561,
     280  =>  3548,
     281  =>  3534,
     282  =>  3521,
     283  =>  3508,
     284  =>  3495,
     285  =>  3482,
     286  =>  3469,
     287  =>  3457,
     288  =>  3444,
     289  =>  3431,
     290  =>  3419,
     291  =>  3407,
     292  =>  3394,
     293  =>  3382,
     294  =>  3370,
     295  =>  3358,
     296  =>  3346,
     297  =>  3334,
     298  =>  3322,
     299  =>  3310,
     300  =>  3299,
     301  =>  3287,
     302  =>  3275,
     303  =>  3264,
     304  =>  3253,
     305  =>  3241,
     306  =>  3230,
     307  =>  3219,
     308  =>  3208,
     309  =>  3197,
     310  =>  3186,
     311  =>  3175,
     312  =>  3164,
     313  =>  3153,
     314  =>  3143,
     315  =>  3132,
     316  =>  3121,
     317  =>  3111,
     318  =>  3100,
     319  =>  3090,
     320  =>  3080,
     321  =>  3069,
     322  =>  3059,
     323  =>  3049,
     324  =>  3039,
     325  =>  3029,
     326  =>  3019,
     327  =>  3009,
     328  =>  2999,
     329  =>  2990,
     330  =>  2980,
     331  =>  2970,
     332  =>  2961,
     333  =>  2951,
     334  =>  2942,
     335  =>  2932,
     336  =>  2923,
     337  =>  2913,
     338  =>  2904,
     339  =>  2895,
     340  =>  2886,
     341  =>  2876,
     342  =>  2867,
     343  =>  2858,
     344  =>  2849,
     345  =>  2840,
     346  =>  2832,
     347  =>  2823,
     348  =>  2814,
     349  =>  2805,
     350  =>  2797,
     351  =>  2788,
     352  =>  2779,
     353  =>  2771,
     354  =>  2762,
     355  =>  2754,
     356  =>  2745,
     357  =>  2737,
     358  =>  2729,
     359  =>  2720,
     360  =>  2712,
     361  =>  2704,
     362  =>  2696,
     363  =>  2688,
     364  =>  2680,
     365  =>  2672,
     366  =>  2664,
     367  =>  2656,
     368  =>  2648,
     369  =>  2640,
     370  =>  2632,
     371  =>  2625,
     372  =>  2617,
     373  =>  2609,
     374  =>  2601,
     375  =>  2594,
     376  =>  2586,
     377  =>  2579,
     378  =>  2571,
     379  =>  2564,
     380  =>  2556,
     381  =>  2549,
     382  =>  2542,
     383  =>  2534,
     384  =>  2527,
     385  =>  2520,
     386  =>  2513,
     387  =>  2505,
     388  =>  2498,
     389  =>  2491,
     390  =>  2484,
     391  =>  2477,
     392  =>  2470,
     393  =>  2463,
     394  =>  2456,
     395  =>  2449,
     396  =>  2442,
     397  =>  2436,
     398  =>  2429,
     399  =>  2422,
     400  =>  2415,
     401  =>  2409,
     402  =>  2402,
     403  =>  2395,
     404  =>  2389,
     405  =>  2382,
     406  =>  2375,
     407  =>  2369,
     408  =>  2362,
     409  =>  2356,
     410  =>  2350,
     411  =>  2343,
     412  =>  2337,
     413  =>  2330,
     414  =>  2324,
     415  =>  2318,
     416  =>  2312,
     417  =>  2305,
     418  =>  2299,
     419  =>  2293,
     420  =>  2287,
     421  =>  2281,
     422  =>  2275,
     423  =>  2269,
     424  =>  2263,
     425  =>  2257,
     426  =>  2251,
     427  =>  2245,
     428  =>  2239,
     429  =>  2233,
     430  =>  2227,
     431  =>  2221,
     432  =>  2215,
     433  =>  2209,
     434  =>  2204,
     435  =>  2198,
     436  =>  2192,
     437  =>  2186,
     438  =>  2181,
     439  =>  2175,
     440  =>  2169,
     441  =>  2164,
     442  =>  2158,
     443  =>  2153,
     444  =>  2147,
     445  =>  2142,
     446  =>  2136,
     447  =>  2131,
     448  =>  2125,
     449  =>  2120,
     450  =>  2114,
     451  =>  2109,
     452  =>  2104,
     453  =>  2098,
     454  =>  2093,
     455  =>  2088,
     456  =>  2082,
     457  =>  2077,
     458  =>  2072,
     459  =>  2067,
     460  =>  2062,
     461  =>  2056,
     462  =>  2051,
     463  =>  2046,
     464  =>  2041,
     465  =>  2036,
     466  =>  2031,
     467  =>  2026,
     468  =>  2021,
     469  =>  2016,
     470  =>  2011,
     471  =>  2006,
     472  =>  2001,
     473  =>  1996,
     474  =>  1991,
     475  =>  1986,
     476  =>  1981,
     477  =>  1977,
     478  =>  1972,
     479  =>  1967,
     480  =>  1962,
     481  =>  1957,
     482  =>  1953,
     483  =>  1948,
     484  =>  1943,
     485  =>  1938,
     486  =>  1934,
     487  =>  1929,
     488  =>  1924,
     489  =>  1920,
     490  =>  1915,
     491  =>  1911,
     492  =>  1906,
     493  =>  1901,
     494  =>  1897,
     495  =>  1892,
     496  =>  1888,
     497  =>  1883,
     498  =>  1879,
     499  =>  1874,
     500  =>  1870,
     501  =>  1866,
     502  =>  1861,
     503  =>  1857,
     504  =>  1852,
     505  =>  1848,
     506  =>  1844,
     507  =>  1839,
     508  =>  1835,
     509  =>  1831,
     510  =>  1826,
     511  =>  1822,
     512  =>  1818,
     513  =>  1814,
     514  =>  1809,
     515  =>  1805,
     516  =>  1801,
     517  =>  1797,
     518  =>  1793,
     519  =>  1788,
     520  =>  1784,
     521  =>  1780,
     522  =>  1776,
     523  =>  1772,
     524  =>  1768,
     525  =>  1764,
     526  =>  1760,
     527  =>  1756,
     528  =>  1752,
     529  =>  1748,
     530  =>  1744,
     531  =>  1740,
     532  =>  1736,
     533  =>  1732,
     534  =>  1728,
     535  =>  1724,
     536  =>  1720,
     537  =>  1716,
     538  =>  1712,
     539  =>  1708,
     540  =>  1704,
     541  =>  1701,
     542  =>  1697,
     543  =>  1693,
     544  =>  1689,
     545  =>  1685,
     546  =>  1681,
     547  =>  1678,
     548  =>  1674,
     549  =>  1670,
     550  =>  1666,
     551  =>  1663,
     552  =>  1659,
     553  =>  1655,
     554  =>  1652,
     555  =>  1648,
     556  =>  1644,
     557  =>  1641,
     558  =>  1637,
     559  =>  1633,
     560  =>  1630,
     561  =>  1626,
     562  =>  1622,
     563  =>  1619,
     564  =>  1615,
     565  =>  1612,
     566  =>  1608,
     567  =>  1605,
     568  =>  1601,
     569  =>  1598,
     570  =>  1594,
     571  =>  1591,
     572  =>  1587,
     573  =>  1584,
     574  =>  1580,
     575  =>  1577,
     576  =>  1573,
     577  =>  1570,
     578  =>  1566,
     579  =>  1563,
     580  =>  1560,
     581  =>  1556,
     582  =>  1553,
     583  =>  1549,
     584  =>  1546,
     585  =>  1543,
     586  =>  1539,
     587  =>  1536,
     588  =>  1533,
     589  =>  1529,
     590  =>  1526,
     591  =>  1523,
     592  =>  1519,
     593  =>  1516,
     594  =>  1513,
     595  =>  1510,
     596  =>  1506,
     597  =>  1503,
     598  =>  1500,
     599  =>  1497,
     600  =>  1494,
     601  =>  1490,
     602  =>  1487,
     603  =>  1484,
     604  =>  1481,
     605  =>  1478,
     606  =>  1475,
     607  =>  1471,
     608  =>  1468,
     609  =>  1465,
     610  =>  1462,
     611  =>  1459,
     612  =>  1456,
     613  =>  1453,
     614  =>  1450,
     615  =>  1447,
     616  =>  1443,
     617  =>  1440,
     618  =>  1437,
     619  =>  1434,
     620  =>  1431,
     621  =>  1428,
     622  =>  1425,
     623  =>  1422,
     624  =>  1419,
     625  =>  1416,
     626  =>  1413,
     627  =>  1410,
     628  =>  1407,
     629  =>  1404,
     630  =>  1401,
     631  =>  1399,
     632  =>  1396,
     633  =>  1393,
     634  =>  1390,
     635  =>  1387,
     636  =>  1384,
     637  =>  1381,
     638  =>  1378,
     639  =>  1375,
     640  =>  1372,
     641  =>  1370,
     642  =>  1367,
     643  =>  1364,
     644  =>  1361,
     645  =>  1358,
     646  =>  1355,
     647  =>  1353,
     648  =>  1350,
     649  =>  1347,
     650  =>  1344,
     651  =>  1341,
     652  =>  1339,
     653  =>  1336,
     654  =>  1333,
     655  =>  1330,
     656  =>  1328,
     657  =>  1325,
     658  =>  1322,
     659  =>  1319,
     660  =>  1317,
     661  =>  1314,
     662  =>  1311,
     663  =>  1309,
     664  =>  1306,
     665  =>  1303,
     666  =>  1301,
     667  =>  1298,
     668  =>  1295,
     669  =>  1293,
     670  =>  1290,
     671  =>  1287,
     672  =>  1285,
     673  =>  1282,
     674  =>  1279,
     675  =>  1277,
     676  =>  1274,
     677  =>  1271,
     678  =>  1269,
     679  =>  1266,
     680  =>  1264,
     681  =>  1261,
     682  =>  1259,
     683  =>  1256,
     684  =>  1253,
     685  =>  1251,
     686  =>  1248,
     687  =>  1246,
     688  =>  1243,
     689  =>  1241,
     690  =>  1238,
     691  =>  1236,
     692  =>  1233,
     693  =>  1231,
     694  =>  1228,
     695  =>  1226,
     696  =>  1223,
     697  =>  1221,
     698  =>  1218,
     699  =>  1216,
     700  =>  1213,
     701  =>  1211,
     702  =>  1208,
     703  =>  1206,
     704  =>  1203,
     705  =>  1201,
     706  =>  1199,
     707  =>  1196,
     708  =>  1194,
     709  =>  1191,
     710  =>  1189,
     711  =>  1187,
     712  =>  1184,
     713  =>  1182,
     714  =>  1179,
     715  =>  1177,
     716  =>  1175,
     717  =>  1172,
     718  =>  1170,
     719  =>  1168,
     720  =>  1165,
     721  =>  1163,
     722  =>  1160,
     723  =>  1158,
     724  =>  1156,
     725  =>  1153,
     726  =>  1151,
     727  =>  1149,
     728  =>  1147,
     729  =>  1144,
     730  =>  1142,
     731  =>  1140,
     732  =>  1137,
     733  =>  1135,
     734  =>  1133,
     735  =>  1131,
     736  =>  1128,
     737  =>  1126,
     738  =>  1124,
     739  =>  1121,
     740  =>  1119,
     741  =>  1117,
     742  =>  1115,
     743  =>  1112,
     744  =>  1110,
     745  =>  1108,
     746  =>  1106,
     747  =>  1104,
     748  =>  1101,
     749  =>  1099,
     750  =>  1097,
     751  =>  1095,
     752  =>  1093,
     753  =>  1090,
     754  =>  1088,
     755  =>  1086,
     756  =>  1084,
     757  =>  1082,
     758  =>  1080,
     759  =>  1077,
     760  =>  1075,
     761  =>  1073,
     762  =>  1071,
     763  =>  1069,
     764  =>  1067,
     765  =>  1065,
     766  =>  1062,
     767  =>  1060,
     768  =>  1058,
     769  =>  1056,
     770  =>  1054,
     771  =>  1052,
     772  =>  1050,
     773  =>  1048,
     774  =>  1046,
     775  =>  1043,
     776  =>  1041,
     777  =>  1039,
     778  =>  1037,
     779  =>  1035,
     780  =>  1033,
     781  =>  1031,
     782  =>  1029,
     783  =>  1027,
     784  =>  1025,
     785  =>  1023,
     786  =>  1021,
     787  =>  1019,
     788  =>  1017,
     789  =>  1015,
     790  =>  1013,
     791  =>  1011,
     792  =>  1009,
     793  =>  1007,
     794  =>  1005,
     795  =>  1003,
     796  =>  1001,
     797  =>   999,
     798  =>   997,
     799  =>   995,
     800  =>   993,
     801  =>   991,
     802  =>   989,
     803  =>   987,
     804  =>   985,
     805  =>   983,
     806  =>   981,
     807  =>   979,
     808  =>   977,
     809  =>   975,
     810  =>   973,
     811  =>   971,
     812  =>   969,
     813  =>   967,
     814  =>   965,
     815  =>   963,
     816  =>   961,
     817  =>   959,
     818  =>   957,
     819  =>   955,
     820  =>   954,
     821  =>   952,
     822  =>   950,
     823  =>   948,
     824  =>   946,
     825  =>   944,
     826  =>   942,
     827  =>   940,
     828  =>   938,
     829  =>   937,
     830  =>   935,
     831  =>   933,
     832  =>   931,
     833  =>   929,
     834  =>   927,
     835  =>   925,
     836  =>   923,
     837  =>   922,
     838  =>   920,
     839  =>   918,
     840  =>   916,
     841  =>   914,
     842  =>   912,
     843  =>   911,
     844  =>   909,
     845  =>   907,
     846  =>   905,
     847  =>   903,
     848  =>   901,
     849  =>   900,
     850  =>   898,
     851  =>   896,
     852  =>   894,
     853  =>   892,
     854  =>   891,
     855  =>   889,
     856  =>   887,
     857  =>   885,
     858  =>   883,
     859  =>   882,
     860  =>   880,
     861  =>   878,
     862  =>   876,
     863  =>   874,
     864  =>   873,
     865  =>   871,
     866  =>   869,
     867  =>   867,
     868  =>   866,
     869  =>   864,
     870  =>   862,
     871  =>   860,
     872  =>   859,
     873  =>   857,
     874  =>   855,
     875  =>   853,
     876  =>   852,
     877  =>   850,
     878  =>   848,
     879  =>   847,
     880  =>   845,
     881  =>   843,
     882  =>   841,
     883  =>   840,
     884  =>   838,
     885  =>   836,
     886  =>   835,
     887  =>   833,
     888  =>   831,
     889  =>   829,
     890  =>   828,
     891  =>   826,
     892  =>   824,
     893  =>   823,
     894  =>   821,
     895  =>   819,
     896  =>   818,
     897  =>   816,
     898  =>   814,
     899  =>   813,
     900  =>   811,
     901  =>   809,
     902  =>   808,
     903  =>   806,
     904  =>   804,
     905  =>   803,
     906  =>   801,
     907  =>   799,
     908  =>   798,
     909  =>   796,
     910  =>   794,
     911  =>   793,
     912  =>   791,
     913  =>   789,
     914  =>   788,
     915  =>   786,
     916  =>   785,
     917  =>   783,
     918  =>   781,
     919  =>   780,
     920  =>   778,
     921  =>   777,
     922  =>   775,
     923  =>   773,
     924  =>   772,
     925  =>   770,
     926  =>   768,
     927  =>   767,
     928  =>   765,
     929  =>   764,
     930  =>   762,
     931  =>   760,
     932  =>   759,
     933  =>   757,
     934  =>   756,
     935  =>   754,
     936  =>   753,
     937  =>   751,
     938  =>   749,
     939  =>   748,
     940  =>   746,
     941  =>   745,
     942  =>   743,
     943  =>   742,
     944  =>   740,
     945  =>   738,
     946  =>   737,
     947  =>   735,
     948  =>   734,
     949  =>   732,
     950  =>   731,
     951  =>   729,
     952  =>   728,
     953  =>   726,
     954  =>   725,
     955  =>   723,
     956  =>   721,
     957  =>   720,
     958  =>   718,
     959  =>   717,
     960  =>   715,
     961  =>   714,
     962  =>   712,
     963  =>   711,
     964  =>   709,
     965  =>   708,
     966  =>   706,
     967  =>   705,
     968  =>   703,
     969  =>   702,
     970  =>   700,
     971  =>   699,
     972  =>   697,
     973  =>   696,
     974  =>   694,
     975  =>   693,
     976  =>   691,
     977  =>   690,
     978  =>   688,
     979  =>   687,
     980  =>   685,
     981  =>   684,
     982  =>   682,
     983  =>   681,
     984  =>   679,
     985  =>   678,
     986  =>   676,
     987  =>   675,
     988  =>   674,
     989  =>   672,
     990  =>   671,
     991  =>   669,
     992  =>   668,
     993  =>   666,
     994  =>   665,
     995  =>   663,
     996  =>   662,
     997  =>   660,
     998  =>   659,
     999  =>   658,
    1000  =>   656,
    1001  =>   655,
    1002  =>   653,
    1003  =>   652,
    1004  =>   650,
    1005  =>   649,
    1006  =>   647,
    1007  =>   646,
    1008  =>   645,
    1009  =>   643,
    1010  =>   642,
    1011  =>   640,
    1012  =>   639,
    1013  =>   637,
    1014  =>   636,
    1015  =>   635,
    1016  =>   633,
    1017  =>   632,
    1018  =>   630,
    1019  =>   629,
    1020  =>   628,
    1021  =>   626,
    1022  =>   625,
    1023  =>   623,
    1024  =>   622,
    1025  =>   621,
    1026  =>   619,
    1027  =>   618,
    1028  =>   616,
    1029  =>   615,
    1030  =>   614,
    1031  =>   612,
    1032  =>   611,
    1033  =>   609,
    1034  =>   608,
    1035  =>   607,
    1036  =>   605,
    1037  =>   604,
    1038  =>   602,
    1039  =>   601,
    1040  =>   600,
    1041  =>   598,
    1042  =>   597,
    1043  =>   596,
    1044  =>   594,
    1045  =>   593,
    1046  =>   591,
    1047  =>   590,
    1048  =>   589,
    1049  =>   587,
    1050  =>   586,
    1051  =>   585,
    1052  =>   583,
    1053  =>   582,
    1054  =>   581,
    1055  =>   579,
    1056  =>   578,
    1057  =>   577,
    1058  =>   575,
    1059  =>   574,
    1060  =>   573,
    1061  =>   571,
    1062  =>   570,
    1063  =>   568,
    1064  =>   567,
    1065  =>   566,
    1066  =>   564,
    1067  =>   563,
    1068  =>   562,
    1069  =>   560,
    1070  =>   559,
    1071  =>   558,
    1072  =>   556,
    1073  =>   555,
    1074  =>   554,
    1075  =>   553,
    1076  =>   551,
    1077  =>   550,
    1078  =>   549,
    1079  =>   547,
    1080  =>   546,
    1081  =>   545,
    1082  =>   543,
    1083  =>   542,
    1084  =>   541,
    1085  =>   539,
    1086  =>   538,
    1087  =>   537,
    1088  =>   535,
    1089  =>   534,
    1090  =>   533,
    1091  =>   532,
    1092  =>   530,
    1093  =>   529,
    1094  =>   528,
    1095  =>   526,
    1096  =>   525,
    1097  =>   524,
    1098  =>   522,
    1099  =>   521,
    1100  =>   520,
    1101  =>   519,
    1102  =>   517,
    1103  =>   516,
    1104  =>   515,
    1105  =>   513,
    1106  =>   512,
    1107  =>   511,
    1108  =>   510,
    1109  =>   508,
    1110  =>   507,
    1111  =>   506,
    1112  =>   505,
    1113  =>   503,
    1114  =>   502,
    1115  =>   501,
    1116  =>   499,
    1117  =>   498,
    1118  =>   497,
    1119  =>   496,
    1120  =>   494,
    1121  =>   493,
    1122  =>   492,
    1123  =>   491,
    1124  =>   489,
    1125  =>   488,
    1126  =>   487,
    1127  =>   486,
    1128  =>   484,
    1129  =>   483,
    1130  =>   482,
    1131  =>   481,
    1132  =>   479,
    1133  =>   478,
    1134  =>   477,
    1135  =>   476,
    1136  =>   474,
    1137  =>   473,
    1138  =>   472,
    1139  =>   471,
    1140  =>   469,
    1141  =>   468,
    1142  =>   467,
    1143  =>   466,
    1144  =>   464,
    1145  =>   463,
    1146  =>   462,
    1147  =>   461,
    1148  =>   459,
    1149  =>   458,
    1150  =>   457,
    1151  =>   456,
    1152  =>   455,
    1153  =>   453,
    1154  =>   452,
    1155  =>   451,
    1156  =>   450,
    1157  =>   448,
    1158  =>   447,
    1159  =>   446,
    1160  =>   445,
    1161  =>   444,
    1162  =>   442,
    1163  =>   441,
    1164  =>   440,
    1165  =>   439,
    1166  =>   438,
    1167  =>   436,
    1168  =>   435,
    1169  =>   434,
    1170  =>   433,
    1171  =>   431,
    1172  =>   430,
    1173  =>   429,
    1174  =>   428,
    1175  =>   427,
    1176  =>   425,
    1177  =>   424,
    1178  =>   423,
    1179  =>   422,
    1180  =>   421,
    1181  =>   419,
    1182  =>   418,
    1183  =>   417,
    1184  =>   416,
    1185  =>   415,
    1186  =>   414,
    1187  =>   412,
    1188  =>   411,
    1189  =>   410,
    1190  =>   409,
    1191  =>   408,
    1192  =>   406,
    1193  =>   405,
    1194  =>   404,
    1195  =>   403,
    1196  =>   402,
    1197  =>   400,
    1198  =>   399,
    1199  =>   398,
    1200  =>   397,
    1201  =>   396,
    1202  =>   395,
    1203  =>   393,
    1204  =>   392,
    1205  =>   391,
    1206  =>   390,
    1207  =>   389,
    1208  =>   388,
    1209  =>   386,
    1210  =>   385,
    1211  =>   384,
    1212  =>   383,
    1213  =>   382,
    1214  =>   381,
    1215  =>   379,
    1216  =>   378,
    1217  =>   377,
    1218  =>   376,
    1219  =>   375,
    1220  =>   374,
    1221  =>   372,
    1222  =>   371,
    1223  =>   370,
    1224  =>   369,
    1225  =>   368,
    1226  =>   367,
    1227  =>   365,
    1228  =>   364,
    1229  =>   363,
    1230  =>   362,
    1231  =>   361,
    1232  =>   360,
    1233  =>   359,
    1234  =>   357,
    1235  =>   356,
    1236  =>   355,
    1237  =>   354,
    1238  =>   353,
    1239  =>   352,
    1240  =>   351,
    1241  =>   349,
    1242  =>   348,
    1243  =>   347,
    1244  =>   346,
    1245  =>   345,
    1246  =>   344,
    1247  =>   343,
    1248  =>   341,
    1249  =>   340,
    1250  =>   339,
    1251  =>   338,
    1252  =>   337,
    1253  =>   336,
    1254  =>   335,
    1255  =>   333,
    1256  =>   332,
    1257  =>   331,
    1258  =>   330,
    1259  =>   329,
    1260  =>   328,
    1261  =>   327,
    1262  =>   326,
    1263  =>   324,
    1264  =>   323,
    1265  =>   322,
    1266  =>   321,
    1267  =>   320,
    1268  =>   319,
    1269  =>   318,
    1270  =>   317,
    1271  =>   315,
    1272  =>   314,
    1273  =>   313,
    1274  =>   312,
    1275  =>   311,
    1276  =>   310,
    1277  =>   309,
    1278  =>   308,
    1279  =>   306,
    1280  =>   305,
    1281  =>   304,
    1282  =>   303,
    1283  =>   302,
    1284  =>   301,
    1285  =>   300,
    1286  =>   299,
    1287  =>   298,
    1288  =>   296,
    1289  =>   295,
    1290  =>   294,
    1291  =>   293,
    1292  =>   292,
    1293  =>   291,
    1294  =>   290,
    1295  =>   289,
    1296  =>   288,
    1297  =>   286,
    1298  =>   285,
    1299  =>   284,
    1300  =>   283,
    1301  =>   282,
    1302  =>   281,
    1303  =>   280,
    1304  =>   279,
    1305  =>   278,
    1306  =>   277,
    1307  =>   275,
    1308  =>   274,
    1309  =>   273,
    1310  =>   272,
    1311  =>   271,
    1312  =>   270,
    1313  =>   269,
    1314  =>   268,
    1315  =>   267,
    1316  =>   266,
    1317  =>   265,
    1318  =>   263,
    1319  =>   262,
    1320  =>   261,
    1321  =>   260,
    1322  =>   259,
    1323  =>   258,
    1324  =>   257,
    1325  =>   256,
    1326  =>   255,
    1327  =>   254,
    1328  =>   253,
    1329  =>   251,
    1330  =>   250,
    1331  =>   249,
    1332  =>   248,
    1333  =>   247,
    1334  =>   246,
    1335  =>   245,
    1336  =>   244,
    1337  =>   243,
    1338  =>   242,
    1339  =>   241,
    1340  =>   240,
    1341  =>   238,
    1342  =>   237,
    1343  =>   236,
    1344  =>   235,
    1345  =>   234,
    1346  =>   233,
    1347  =>   232,
    1348  =>   231,
    1349  =>   230,
    1350  =>   229,
    1351  =>   228,
    1352  =>   227,
    1353  =>   226,
    1354  =>   224,
    1355  =>   223,
    1356  =>   222,
    1357  =>   221,
    1358  =>   220,
    1359  =>   219,
    1360  =>   218,
    1361  =>   217,
    1362  =>   216,
    1363  =>   215,
    1364  =>   214,
    1365  =>   213,
    1366  =>   212,
    1367  =>   211,
    1368  =>   209,
    1369  =>   208,
    1370  =>   207,
    1371  =>   206,
    1372  =>   205,
    1373  =>   204,
    1374  =>   203,
    1375  =>   202,
    1376  =>   201,
    1377  =>   200,
    1378  =>   199,
    1379  =>   198,
    1380  =>   197,
    1381  =>   196,
    1382  =>   195,
    1383  =>   194,
    1384  =>   192,
    1385  =>   191,
    1386  =>   190,
    1387  =>   189,
    1388  =>   188,
    1389  =>   187,
    1390  =>   186,
    1391  =>   185,
    1392  =>   184,
    1393  =>   183,
    1394  =>   182,
    1395  =>   181,
    1396  =>   180,
    1397  =>   179,
    1398  =>   178,
    1399  =>   177,
    1400  =>   176,
    1401  =>   175,
    1402  =>   173,
    1403  =>   172,
    1404  =>   171,
    1405  =>   170,
    1406  =>   169,
    1407  =>   168,
    1408  =>   167,
    1409  =>   166,
    1410  =>   165,
    1411  =>   164,
    1412  =>   163,
    1413  =>   162,
    1414  =>   161,
    1415  =>   160,
    1416  =>   159,
    1417  =>   158,
    1418  =>   157,
    1419  =>   156,
    1420  =>   155,
    1421  =>   154,
    1422  =>   152,
    1423  =>   151,
    1424  =>   150,
    1425  =>   149,
    1426  =>   148,
    1427  =>   147,
    1428  =>   146,
    1429  =>   145,
    1430  =>   144,
    1431  =>   143,
    1432  =>   142,
    1433  =>   141,
    1434  =>   140,
    1435  =>   139,
    1436  =>   138,
    1437  =>   137,
    1438  =>   136,
    1439  =>   135,
    1440  =>   134,
    1441  =>   133,
    1442  =>   132,
    1443  =>   131,
    1444  =>   129,
    1445  =>   128,
    1446  =>   127,
    1447  =>   126,
    1448  =>   125,
    1449  =>   124,
    1450  =>   123,
    1451  =>   122,
    1452  =>   121,
    1453  =>   120,
    1454  =>   119,
    1455  =>   118,
    1456  =>   117,
    1457  =>   116,
    1458  =>   115,
    1459  =>   114,
    1460  =>   113,
    1461  =>   112,
    1462  =>   111,
    1463  =>   110,
    1464  =>   109,
    1465  =>   108,
    1466  =>   107,
    1467  =>   106,
    1468  =>   105,
    1469  =>   104,
    1470  =>   103,
    1471  =>   101,
    1472  =>   100,
    1473  =>    99,
    1474  =>    98,
    1475  =>    97,
    1476  =>    96,
    1477  =>    95,
    1478  =>    94,
    1479  =>    93,
    1480  =>    92,
    1481  =>    91,
    1482  =>    90,
    1483  =>    89,
    1484  =>    88,
    1485  =>    87,
    1486  =>    86,
    1487  =>    85,
    1488  =>    84,
    1489  =>    83,
    1490  =>    82,
    1491  =>    81,
    1492  =>    80,
    1493  =>    79,
    1494  =>    78,
    1495  =>    77,
    1496  =>    76,
    1497  =>    75,
    1498  =>    74,
    1499  =>    73,
    1500  =>    72,
    1501  =>    71,
    1502  =>    70,
    1503  =>    69,
    1504  =>    67,
    1505  =>    66,
    1506  =>    65,
    1507  =>    64,
    1508  =>    63,
    1509  =>    62,
    1510  =>    61,
    1511  =>    60,
    1512  =>    59,
    1513  =>    58,
    1514  =>    57,
    1515  =>    56,
    1516  =>    55,
    1517  =>    54,
    1518  =>    53,
    1519  =>    52,
    1520  =>    51,
    1521  =>    50,
    1522  =>    49,
    1523  =>    48,
    1524  =>    47,
    1525  =>    46,
    1526  =>    45,
    1527  =>    44,
    1528  =>    43,
    1529  =>    42,
    1530  =>    41,
    1531  =>    40,
    1532  =>    39,
    1533  =>    38,
    1534  =>    37,
    1535  =>    36,
    1536  =>    35,
    1537  =>    34,
    1538  =>    33,
    1539  =>    32,
    1540  =>    31,
    1541  =>    29,
    1542  =>    28,
    1543  =>    27,
    1544  =>    26,
    1545  =>    25,
    1546  =>    24,
    1547  =>    23,
    1548  =>    22,
    1549  =>    21,
    1550  =>    20,
    1551  =>    19,
    1552  =>    18,
    1553  =>    17,
    1554  =>    16,
    1555  =>    15,
    1556  =>    14,
    1557  =>    13,
    1558  =>    12,
    1559  =>    11,
    1560  =>    10,
    1561  =>     9,
    1562  =>     8,
    1563  =>     7,
    1564  =>     6,
    1565  =>     5,
    1566  =>     4,
    1567  =>     3,
    1568  =>     2
  );

 end package roi_tan;
