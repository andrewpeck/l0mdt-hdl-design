--------------------------------------------------------------------------------
--  UMass , Physics Department
--  Guillermo Loustau de Linares
--  gloustau@cern.ch
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger
--  Module: Trigonometrics functions
--  Description: 
--      Readers for: tan & arctan
--            
--------------------------------------------------------------------------------
--  Revisions:
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package roi_trig_functions is
  
  
  
end package roi_trig_functions;

package body roi_trig_functions is
  
  
  
end package body roi_trig_functions;