class Rand40;
   rand bit l1a_req;

   //constraint src {
   //   l1a_req dist { 1'b0 := 49, 1'b1 := 1 };
   //}
   
endclass // Transaction
