--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: angle to tube number offset
--  Multiplier: 1 
--  slope are defined with angle relative to beam line
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library heg_roi_lib;
use heg_roi_lib.roi_types_pkg.all;

package roi_lut_BILA3_slope is

  -- add length of constant array
  constant ROM_BILA3_ANGLE_MAX_SIZE : integer := 2048;

-- VHDL2008  -- constant ROI_BILA3_SLOPE_MEM : roi_mbar_lut_t(ROM_BILA3_SLOPE_MAX_SIZE - 1 downto 0)(0 to 5) := (
  constant ROI_BILA3_ANGLE_MEM : roi_mbar_lut_large_t(ROM_BILA3_ANGLE_MAX_SIZE - 1 downto 0) := (
   2047 downto  366 => ( ( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5) ), -- from 89.10482629 to 85 degree 
    365 downto  119 => ( ( -6,  4),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -4,  6) ), -- from 85 to 75 degree 
    118 downto   69 => ( ( -7,  3),( -6,  4),( -6,  4),( -6,  4),( -4,  6),( -4,  6),( -4,  6),( -3,  7) ), -- from 75 to 65 degree 
     68 downto   46 => ( ( -8,  2),( -8,  2),( -7,  3),( -6,  4),( -4,  6),( -3,  7),( -2,  8),( -2,  8) ), -- from 65 to 55 degree 
     45 downto   38 => ( ( -9,  1),( -9,  1),( -8,  2),( -7,  3),( -3,  7),( -2,  8),( -1,  9),( -1,  9) ), -- from 55 to 50 degree 
     37 downto   32 => ( (-10,  0),( -9,  1),( -8,  2),( -8,  2),( -2,  8),( -2,  8),( -1,  9),(  0, 10) ), -- from 50 to 45 degree 
     31 downto   27 => ( (-11, -1),(-10,  0),( -9,  1),( -8,  2),( -2,  8),( -1,  9),(  0, 10),(  1, 11) ), -- from 45 to 40 degree 
     26 downto   22 => ( (-13, -3),(-11, -1),(-10,  0),( -9,  1),( -1,  9),(  0, 10),(  1, 11),(  3, 13) ), -- from 40 to 35 degree 
     21 downto   18 => ( (-14, -4),(-13, -3),(-11, -1),(-10,  0),(  0, 10),(  1, 11),(  3, 13),(  4, 14) ), -- from 35 to 30 degree 
     17 downto   15 => ( (-17, -7),(-15, -5),(-13, -3),(-11, -1),(  1, 11),(  3, 13),(  5, 15),(  7, 17) ), -- from 30 to 25 degree 
     14 downto   12 => ( (-20,-10),(-17, -7),(-15, -5),(-13, -3),(  3, 13),(  5, 15),(  7, 17),( 10, 20) ), -- from 25 to 20 degree 
     11 downto    9 => ( (-25,-15),(-21,-11),(-18, -8),(-15, -5),(  5, 15),(  8, 18),( 11, 21),( 15, 25) ), -- from 20 to 15 degree 
      8 downto    6 => ( (-33,-23),(-29,-19),(-24,-14),(-20,-10),( 10, 20),( 14, 24),( 19, 29),( 23, 33) ), -- from 15 to 10 degree 
      5 downto    0 => ( (-53,-43),(-45,-35),(-37,-27),(-30,-20),( 20, 30),( 27, 37),( 35, 45),( 43, 53) )  -- from 10 to 5 degree 
  );

 end package roi_lut_BILA3_slope;

