--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: angle to tube number offset
--  Multiplier: 1 
--  slope are defined with angle relative to beam line
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library heg_roi_lib;
use heg_roi_lib.roi_types_pkg.all;

package roi_lut_BMLA3_slope is

  -- add length of constant array
  constant ROM_BMLA3_ANGLE_MAX_SIZE : integer := 2048;

-- VHDL2008  -- constant ROI_BMLA3_SLOPE_MEM : roi_mbar_lut_t(ROM_BMLA3_SLOPE_MAX_SIZE - 1 downto 0)(0 to 5) := (
  constant ROI_BMLA3_ANGLE_MEM : roi_mbar_lut_small_t(ROM_BMLA3_ANGLE_MAX_SIZE - 1 downto 0) := (
    2047 downto 1921 => ( ( -2,  8),( -3,  7),( -3,  7),( -7,  3),( -7,  3),( -8,  2) ), -- from 117.28 to 110 degree 
    1920 downto 1834 => ( ( -3,  7),( -3,  7),( -4,  6),( -6,  4),( -7,  3),( -7,  3) ), -- from 110 to 105 degree 
    1833 downto 1746 => ( ( -4,  6),( -4,  6),( -4,  6),( -6,  4),( -6,  4),( -6,  4) ), -- from 105 to 100 degree 
    1745 downto 1659 => ( ( -4,  6),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -6,  4) ), -- from 100 to 95 degree 
    1658 downto 1485 => ( ( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5),( -5,  5) ), -- from 95 to 85 degree 
    1484 downto 1310 => ( ( -6,  4),( -6,  4),( -6,  4),( -4,  6),( -4,  6),( -4,  6) ), -- from 85 to 75 degree 
    1309 downto 1135 => ( ( -7,  3),( -7,  3),( -7,  3),( -3,  7),( -3,  7),( -3,  7) ), -- from 75 to 65 degree 
    1134 downto  961 => ( ( -9,  1),( -8,  2),( -8,  2),( -2,  8),( -2,  8),( -1,  9) ), -- from 65 to 55 degree 
     960 downto  874 => ( (-10,  0),(-10,  0),( -9,  1),( -1,  9),(  0, 10),(  0, 10) ), -- from 55 to 50 degree 
     873 downto  786 => ( (-12, -2),(-11, -1),(-10,  0),(  0, 10),(  1, 11),(  2, 12) ), -- from 50 to 45 degree 
     785 downto  699 => ( (-13, -3),(-12, -2),(-11, -1),(  1, 11),(  2, 12),(  3, 13) ), -- from 45 to 40 degree 
     698 downto  612 => ( (-15, -5),(-13, -3),(-12, -2),(  2, 12),(  3, 13),(  5, 15) ), -- from 40 to 35 degree 
     611 downto  525 => ( (-17, -7),(-15, -5),(-14, -4),(  4, 14),(  5, 15),(  7, 17) ), -- from 35 to 30 degree 
     524 downto  437 => ( (-19, -9),(-18, -8),(-16, -6),(  6, 16),(  8, 18),(  9, 19) ), -- from 30 to 25 degree 
     436 downto  350 => ( (-23,-13),(-21,-11),(-18, -8),(  8, 18),( 11, 21),( 13, 23) ), -- from 25 to 20 degree 
     349 downto  263 => ( (-29,-19),(-26,-16),(-23,-13),( 13, 23),( 16, 26),( 19, 29) ), -- from 20 to 15 degree 
     262 downto  176 => ( (-40,-30),(-35,-25),(-31,-21),( 21, 31),( 25, 35),( 30, 40) ), -- from 15 to 10 degree 
     175 downto    0 => ( (-64,-54),(-56,-46),(-48,-38),( 38, 48),( 46, 56),( 54, 64) )  -- from 10 to 5 degree 
  );

 end package roi_lut_BMLA3_slope;

