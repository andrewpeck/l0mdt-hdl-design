library ieee;
use ieee.std_logic_1164.all;
package c2cslave_pkg is
  component c2cSlave is
  port (
    clk50Mhz : in STD_LOGIC;
    reset_n : in STD_LOGIC;
    AXI_CLK : in STD_LOGIC;
    AXI_RST_N : out std_logic;
    K_C2CLINK_aurora_do_cc : out STD_LOGIC;
    K_C2CLINK_axi_c2c_config_error_out : out STD_LOGIC;
    K_C2CLINK_axi_c2c_link_status_out : out STD_LOGIC;
    K_C2CLINK_axi_c2c_multi_bit_error_out : out STD_LOGIC;
    K_C2CLINK_PHY_power_down : in STD_LOGIC;
    K_C2CLINK_PHY_gt_pll_lock : out STD_LOGIC;
    K_C2CLINK_PHY_hard_err : out STD_LOGIC;
    K_C2CLINK_PHY_soft_err : out STD_LOGIC;
    K_C2CLINK_PHY_lane_up : out std_logic;
    K_C2CLINK_PHY_mmcm_not_locked_out : out STD_LOGIC;
    K_C2CLINK_PHY_link_reset_out : out STD_LOGIC;
    KINTEX_SYS_MGMT_alarm : out STD_LOGIC;
    KINTEX_SYS_MGMT_vccint_alarm : out STD_LOGIC;
    KINTEX_SYS_MGMT_vccaux_alarm : out STD_LOGIC;
    KINTEX_SYS_MGMT_overtemp_alarm : out STD_LOGIC;
    clk40 : in STD_LOGIC;
    FW_INFO_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    FW_INFO_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    FW_INFO_awvalid : out STD_LOGIC;
    FW_INFO_awready : in STD_LOGIC;
    FW_INFO_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    FW_INFO_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    FW_INFO_wvalid : out STD_LOGIC;
    FW_INFO_wready : in STD_LOGIC;
    FW_INFO_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    FW_INFO_bvalid : in STD_LOGIC;
    FW_INFO_bready : out STD_LOGIC;
    FW_INFO_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    FW_INFO_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    FW_INFO_arvalid : out STD_LOGIC;
    FW_INFO_arready : in STD_LOGIC;
    FW_INFO_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    FW_INFO_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    FW_INFO_rvalid : in STD_LOGIC;
    FW_INFO_rready : out STD_LOGIC;
    HAL_CORE_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_CORE_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    HAL_CORE_awvalid : out STD_LOGIC;
    HAL_CORE_awready : in STD_LOGIC;
    HAL_CORE_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_CORE_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    HAL_CORE_wvalid : out STD_LOGIC;
    HAL_CORE_wready : in STD_LOGIC;
    HAL_CORE_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    HAL_CORE_bvalid : in STD_LOGIC;
    HAL_CORE_bready : out STD_LOGIC;
    HAL_CORE_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_CORE_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    HAL_CORE_arvalid : out STD_LOGIC;
    HAL_CORE_arready : in STD_LOGIC;
    HAL_CORE_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_CORE_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    HAL_CORE_rvalid : in STD_LOGIC;
    HAL_CORE_rready : out STD_LOGIC;
    UCM_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    UCM_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    UCM_awvalid : out STD_LOGIC;
    UCM_awready : in STD_LOGIC;
    UCM_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    UCM_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    UCM_wvalid : out STD_LOGIC;
    UCM_wready : in STD_LOGIC;
    UCM_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    UCM_bvalid : in STD_LOGIC;
    UCM_bready : out STD_LOGIC;
    UCM_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    UCM_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    UCM_arvalid : out STD_LOGIC;
    UCM_arready : in STD_LOGIC;
    UCM_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    UCM_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    UCM_rvalid : in STD_LOGIC;
    UCM_rready : out STD_LOGIC;
    TAR_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    TAR_awvalid : out STD_LOGIC;
    TAR_awready : in STD_LOGIC;
    TAR_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    TAR_wvalid : out STD_LOGIC;
    TAR_wready : in STD_LOGIC;
    TAR_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    TAR_bvalid : in STD_LOGIC;
    TAR_bready : out STD_LOGIC;
    TAR_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    TAR_arvalid : out STD_LOGIC;
    TAR_arready : in STD_LOGIC;
    TAR_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    TAR_rvalid : in STD_LOGIC;
    TAR_rready : out STD_LOGIC;
    MPL_SPY_PORT_A_addr : out STD_LOGIC_VECTOR ( 14 downto 0 );
    MPL_SPY_PORT_A_clk : out STD_LOGIC;
    MPL_SPY_PORT_A_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_SPY_PORT_A_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_SPY_PORT_A_en : out STD_LOGIC;
    MPL_SPY_PORT_A_rst : out STD_LOGIC;
    MPL_SPY_PORT_A_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    TAR_SPY_PORT_A_addr : out STD_LOGIC_VECTOR ( 15 downto 0 );
    TAR_SPY_PORT_A_clk : out STD_LOGIC;
    TAR_SPY_PORT_A_din : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_SPY_PORT_A_dout : in STD_LOGIC_VECTOR ( 31 downto 0 );
    TAR_SPY_PORT_A_en : out STD_LOGIC;
    TAR_SPY_PORT_A_rst : out STD_LOGIC;
    TAR_SPY_PORT_A_we : out STD_LOGIC_VECTOR ( 3 downto 0 );
    K_C2CLINK_PHY_Tx_txn : out std_logic;
    K_C2CLINK_PHY_Tx_txp : out std_logic;
    K_C2CLINK_PHY_Rx_rxn : in std_logic;
    K_C2CLINK_PHY_Rx_rxp : in std_logic;
    HAL_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    HAL_awvalid : out STD_LOGIC;
    HAL_awready : in STD_LOGIC;
    HAL_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    HAL_wvalid : out STD_LOGIC;
    HAL_wready : in STD_LOGIC;
    HAL_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    HAL_bvalid : in STD_LOGIC;
    HAL_bready : out STD_LOGIC;
    HAL_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    HAL_arvalid : out STD_LOGIC;
    HAL_arready : in STD_LOGIC;
    HAL_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    HAL_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    HAL_rvalid : in STD_LOGIC;
    HAL_rready : out STD_LOGIC;
    K_C2CLINK_PHY_refclk_clk_n : in STD_LOGIC;
    K_C2CLINK_PHY_refclk_clk_p : in STD_LOGIC;
    TF_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TF_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    TF_awvalid : out STD_LOGIC;
    TF_awready : in STD_LOGIC;
    TF_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TF_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    TF_wvalid : out STD_LOGIC;
    TF_wready : in STD_LOGIC;
    TF_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    TF_bvalid : in STD_LOGIC;
    TF_bready : out STD_LOGIC;
    TF_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    TF_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    TF_arvalid : out STD_LOGIC;
    TF_arready : in STD_LOGIC;
    TF_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    TF_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    TF_rvalid : in STD_LOGIC;
    TF_rready : out STD_LOGIC;
    MTC_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MTC_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    MTC_awvalid : out STD_LOGIC;
    MTC_awready : in STD_LOGIC;
    MTC_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MTC_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    MTC_wvalid : out STD_LOGIC;
    MTC_wready : in STD_LOGIC;
    MTC_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    MTC_bvalid : in STD_LOGIC;
    MTC_bready : out STD_LOGIC;
    MTC_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MTC_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    MTC_arvalid : out STD_LOGIC;
    MTC_arready : in STD_LOGIC;
    MTC_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    MTC_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    MTC_rvalid : in STD_LOGIC;
    MTC_rready : out STD_LOGIC;
    DAQ_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    DAQ_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    DAQ_awvalid : out STD_LOGIC;
    DAQ_awready : in STD_LOGIC;
    DAQ_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    DAQ_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    DAQ_wvalid : out STD_LOGIC;
    DAQ_wready : in STD_LOGIC;
    DAQ_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    DAQ_bvalid : in STD_LOGIC;
    DAQ_bready : out STD_LOGIC;
    DAQ_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    DAQ_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    DAQ_arvalid : out STD_LOGIC;
    DAQ_arready : in STD_LOGIC;
    DAQ_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    DAQ_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    DAQ_rvalid : in STD_LOGIC;
    DAQ_rready : out STD_LOGIC;
    H2S_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    H2S_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    H2S_awvalid : out STD_LOGIC;
    H2S_awready : in STD_LOGIC;
    H2S_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    H2S_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    H2S_wvalid : out STD_LOGIC;
    H2S_wready : in STD_LOGIC;
    H2S_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    H2S_bvalid : in STD_LOGIC;
    H2S_bready : out STD_LOGIC;
    H2S_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    H2S_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    H2S_arvalid : out STD_LOGIC;
    H2S_arready : in STD_LOGIC;
    H2S_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    H2S_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    H2S_rvalid : in STD_LOGIC;
    H2S_rready : out STD_LOGIC;
    MPL_awaddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_awprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    MPL_awvalid : out STD_LOGIC;
    MPL_awready : in STD_LOGIC;
    MPL_wdata : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_wstrb : out STD_LOGIC_VECTOR ( 3 downto 0 );
    MPL_wvalid : out STD_LOGIC;
    MPL_wready : in STD_LOGIC;
    MPL_bresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    MPL_bvalid : in STD_LOGIC;
    MPL_bready : out STD_LOGIC;
    MPL_araddr : out STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_arprot : out STD_LOGIC_VECTOR ( 2 downto 0 );
    MPL_arvalid : out STD_LOGIC;
    MPL_arready : in STD_LOGIC;
    MPL_rdata : in STD_LOGIC_VECTOR ( 31 downto 0 );
    MPL_rresp : in STD_LOGIC_VECTOR ( 1 downto 0 );
    MPL_rvalid : in STD_LOGIC;
    MPL_rready : out STD_LOGIC
  );
  end component c2cSlave;
end package c2cslave_pkg;
