--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: slope to angle (mrad) 
--  Multiplier: 2048 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package roi_atan is

    -- add length of constant array
    constant ROM_ATAN_MAX_SIZE : integer := 732388;
    type roi_atan_lut_t is array (integer range <>) of integer;


    constant ROI_ATAN_MEM : roi_atan_lut_t(0 to ROM_ATAN_MAX_SIZE - 1) := (

        0 to     0 =>    0,
        1 to     2 =>    1,
        3 to     4 =>    2,
        5 to     6 =>    3,
        7 to     8 =>    4,
        9 to    10 =>    5,
       11 to    12 =>    6,
       13 to    14 =>    7,
       15 to    16 =>    8,
       17 to    18 =>    9,
       19 to    21 =>   10,
       22 to    23 =>   11,
       24 to    25 =>   12,
       26 to    27 =>   13,
       28 to    29 =>   14,
       30 to    31 =>   15,
       32 to    33 =>   16,
       34 to    35 =>   17,
       36 to    37 =>   18,
       38 to    39 =>   19,
       40 to    41 =>   20,
       42 to    43 =>   21,
       44 to    45 =>   22,
       46 to    47 =>   23,
       48 to    49 =>   24,
       50 to    51 =>   25,
       52 to    53 =>   26,
       54 to    55 =>   27,
       56 to    57 =>   28,
       58 to    59 =>   29,
       60 to    61 =>   30,
       62 to    64 =>   31,
       65 to    66 =>   32,
       67 to    68 =>   33,
       69 to    70 =>   34,
       71 to    72 =>   35,
       73 to    74 =>   36,
       75 to    76 =>   37,
       77 to    78 =>   38,
       79 to    80 =>   39,
       81 to    82 =>   40,
       83 to    84 =>   41,
       85 to    86 =>   42,
       87 to    88 =>   43,
       89 to    90 =>   44,
       91 to    92 =>   45,
       93 to    94 =>   46,
       95 to    96 =>   47,
       97 to    98 =>   48,
       99 to   100 =>   49,
      101 to   103 =>   50,
      104 to   105 =>   51,
      106 to   107 =>   52,
      108 to   109 =>   53,
      110 to   111 =>   54,
      112 to   113 =>   55,
      114 to   115 =>   56,
      116 to   117 =>   57,
      118 to   119 =>   58,
      120 to   121 =>   59,
      122 to   123 =>   60,
      124 to   125 =>   61,
      126 to   127 =>   62,
      128 to   129 =>   63,
      130 to   131 =>   64,
      132 to   133 =>   65,
      134 to   135 =>   66,
      136 to   137 =>   67,
      138 to   140 =>   68,
      141 to   142 =>   69,
      143 to   144 =>   70,
      145 to   146 =>   71,
      147 to   148 =>   72,
      149 to   150 =>   73,
      151 to   152 =>   74,
      153 to   154 =>   75,
      155 to   156 =>   76,
      157 to   158 =>   77,
      159 to   160 =>   78,
      161 to   162 =>   79,
      163 to   164 =>   80,
      165 to   166 =>   81,
      167 to   168 =>   82,
      169 to   170 =>   83,
      171 to   172 =>   84,
      173 to   175 =>   85,
      176 to   177 =>   86,
      178 to   179 =>   87,
      180 to   181 =>   88,
      182 to   183 =>   89,
      184 to   185 =>   90,
      186 to   187 =>   91,
      188 to   189 =>   92,
      190 to   191 =>   93,
      192 to   193 =>   94,
      194 to   195 =>   95,
      196 to   197 =>   96,
      198 to   199 =>   97,
      200 to   201 =>   98,
      202 to   203 =>   99,
      204 to   206 =>  100,
      207 to   208 =>  101,
      209 to   210 =>  102,
      211 to   212 =>  103,
      213 to   214 =>  104,
      215 to   216 =>  105,
      217 to   218 =>  106,
      219 to   220 =>  107,
      221 to   222 =>  108,
      223 to   224 =>  109,
      225 to   226 =>  110,
      227 to   228 =>  111,
      229 to   230 =>  112,
      231 to   232 =>  113,
      233 to   235 =>  114,
      236 to   237 =>  115,
      238 to   239 =>  116,
      240 to   241 =>  117,
      242 to   243 =>  118,
      244 to   245 =>  119,
      246 to   247 =>  120,
      248 to   249 =>  121,
      250 to   251 =>  122,
      252 to   253 =>  123,
      254 to   255 =>  124,
      256 to   257 =>  125,
      258 to   259 =>  126,
      260 to   262 =>  127,
      263 to   264 =>  128,
      265 to   266 =>  129,
      267 to   268 =>  130,
      269 to   270 =>  131,
      271 to   272 =>  132,
      273 to   274 =>  133,
      275 to   276 =>  134,
      277 to   278 =>  135,
      279 to   280 =>  136,
      281 to   282 =>  137,
      283 to   284 =>  138,
      285 to   287 =>  139,
      288 to   289 =>  140,
      290 to   291 =>  141,
      292 to   293 =>  142,
      294 to   295 =>  143,
      296 to   297 =>  144,
      298 to   299 =>  145,
      300 to   301 =>  146,
      302 to   303 =>  147,
      304 to   305 =>  148,
      306 to   307 =>  149,
      308 to   310 =>  150,
      311 to   312 =>  151,
      313 to   314 =>  152,
      315 to   316 =>  153,
      317 to   318 =>  154,
      319 to   320 =>  155,
      321 to   322 =>  156,
      323 to   324 =>  157,
      325 to   326 =>  158,
      327 to   328 =>  159,
      329 to   331 =>  160,
      332 to   333 =>  161,
      334 to   335 =>  162,
      336 to   337 =>  163,
      338 to   339 =>  164,
      340 to   341 =>  165,
      342 to   343 =>  166,
      344 to   345 =>  167,
      346 to   347 =>  168,
      348 to   349 =>  169,
      350 to   352 =>  170,
      353 to   354 =>  171,
      355 to   356 =>  172,
      357 to   358 =>  173,
      359 to   360 =>  174,
      361 to   362 =>  175,
      363 to   364 =>  176,
      365 to   366 =>  177,
      367 to   369 =>  178,
      370 to   371 =>  179,
      372 to   373 =>  180,
      374 to   375 =>  181,
      376 to   377 =>  182,
      378 to   379 =>  183,
      380 to   381 =>  184,
      382 to   383 =>  185,
      384 to   385 =>  186,
      386 to   388 =>  187,
      389 to   390 =>  188,
      391 to   392 =>  189,
      393 to   394 =>  190,
      395 to   396 =>  191,
      397 to   398 =>  192,
      399 to   400 =>  193,
      401 to   402 =>  194,
      403 to   405 =>  195,
      406 to   407 =>  196,
      408 to   409 =>  197,
      410 to   411 =>  198,
      412 to   413 =>  199,
      414 to   415 =>  200,
      416 to   417 =>  201,
      418 to   419 =>  202,
      420 to   422 =>  203,
      423 to   424 =>  204,
      425 to   426 =>  205,
      427 to   428 =>  206,
      429 to   430 =>  207,
      431 to   432 =>  208,
      433 to   434 =>  209,
      435 to   437 =>  210,
      438 to   439 =>  211,
      440 to   441 =>  212,
      442 to   443 =>  213,
      444 to   445 =>  214,
      446 to   447 =>  215,
      448 to   449 =>  216,
      450 to   452 =>  217,
      453 to   454 =>  218,
      455 to   456 =>  219,
      457 to   458 =>  220,
      459 to   460 =>  221,
      461 to   462 =>  222,
      463 to   465 =>  223,
      466 to   467 =>  224,
      468 to   469 =>  225,
      470 to   471 =>  226,
      472 to   473 =>  227,
      474 to   475 =>  228,
      476 to   477 =>  229,
      478 to   480 =>  230,
      481 to   482 =>  231,
      483 to   484 =>  232,
      485 to   486 =>  233,
      487 to   488 =>  234,
      489 to   490 =>  235,
      491 to   493 =>  236,
      494 to   495 =>  237,
      496 to   497 =>  238,
      498 to   499 =>  239,
      500 to   501 =>  240,
      502 to   503 =>  241,
      504 to   506 =>  242,
      507 to   508 =>  243,
      509 to   510 =>  244,
      511 to   512 =>  245,
      513 to   514 =>  246,
      515 to   516 =>  247,
      517 to   519 =>  248,
      520 to   521 =>  249,
      522 to   523 =>  250,
      524 to   525 =>  251,
      526 to   527 =>  252,
      528 to   530 =>  253,
      531 to   532 =>  254,
      533 to   534 =>  255,
      535 to   536 =>  256,
      537 to   538 =>  257,
      539 to   541 =>  258,
      542 to   543 =>  259,
      544 to   545 =>  260,
      546 to   547 =>  261,
      548 to   549 =>  262,
      550 to   551 =>  263,
      552 to   554 =>  264,
      555 to   556 =>  265,
      557 to   558 =>  266,
      559 to   560 =>  267,
      561 to   562 =>  268,
      563 to   565 =>  269,
      566 to   567 =>  270,
      568 to   569 =>  271,
      570 to   571 =>  272,
      572 to   574 =>  273,
      575 to   576 =>  274,
      577 to   578 =>  275,
      579 to   580 =>  276,
      581 to   582 =>  277,
      583 to   585 =>  278,
      586 to   587 =>  279,
      588 to   589 =>  280,
      590 to   591 =>  281,
      592 to   593 =>  282,
      594 to   596 =>  283,
      597 to   598 =>  284,
      599 to   600 =>  285,
      601 to   602 =>  286,
      603 to   605 =>  287,
      606 to   607 =>  288,
      608 to   609 =>  289,
      610 to   611 =>  290,
      612 to   613 =>  291,
      614 to   616 =>  292,
      617 to   618 =>  293,
      619 to   620 =>  294,
      621 to   622 =>  295,
      623 to   625 =>  296,
      626 to   627 =>  297,
      628 to   629 =>  298,
      630 to   631 =>  299,
      632 to   634 =>  300,
      635 to   636 =>  301,
      637 to   638 =>  302,
      639 to   640 =>  303,
      641 to   643 =>  304,
      644 to   645 =>  305,
      646 to   647 =>  306,
      648 to   649 =>  307,
      650 to   652 =>  308,
      653 to   654 =>  309,
      655 to   656 =>  310,
      657 to   658 =>  311,
      659 to   661 =>  312,
      662 to   663 =>  313,
      664 to   665 =>  314,
      666 to   667 =>  315,
      668 to   670 =>  316,
      671 to   672 =>  317,
      673 to   674 =>  318,
      675 to   677 =>  319,
      678 to   679 =>  320,
      680 to   681 =>  321,
      682 to   683 =>  322,
      684 to   686 =>  323,
      687 to   688 =>  324,
      689 to   690 =>  325,
      691 to   692 =>  326,
      693 to   695 =>  327,
      696 to   697 =>  328,
      698 to   699 =>  329,
      700 to   702 =>  330,
      703 to   704 =>  331,
      705 to   706 =>  332,
      707 to   709 =>  333,
      710 to   711 =>  334,
      712 to   713 =>  335,
      714 to   715 =>  336,
      716 to   718 =>  337,
      719 to   720 =>  338,
      721 to   722 =>  339,
      723 to   725 =>  340,
      726 to   727 =>  341,
      728 to   729 =>  342,
      730 to   732 =>  343,
      733 to   734 =>  344,
      735 to   736 =>  345,
      737 to   738 =>  346,
      739 to   741 =>  347,
      742 to   743 =>  348,
      744 to   745 =>  349,
      746 to   748 =>  350,
      749 to   750 =>  351,
      751 to   752 =>  352,
      753 to   755 =>  353,
      756 to   757 =>  354,
      758 to   759 =>  355,
      760 to   762 =>  356,
      763 to   764 =>  357,
      765 to   766 =>  358,
      767 to   769 =>  359,
      770 to   771 =>  360,
      772 to   773 =>  361,
      774 to   776 =>  362,
      777 to   778 =>  363,
      779 to   780 =>  364,
      781 to   783 =>  365,
      784 to   785 =>  366,
      786 to   787 =>  367,
      788 to   790 =>  368,
      791 to   792 =>  369,
      793 to   795 =>  370,
      796 to   797 =>  371,
      798 to   799 =>  372,
      800 to   802 =>  373,
      803 to   804 =>  374,
      805 to   806 =>  375,
      807 to   809 =>  376,
      810 to   811 =>  377,
      812 to   813 =>  378,
      814 to   816 =>  379,
      817 to   818 =>  380,
      819 to   821 =>  381,
      822 to   823 =>  382,
      824 to   825 =>  383,
      826 to   828 =>  384,
      829 to   830 =>  385,
      831 to   832 =>  386,
      833 to   835 =>  387,
      836 to   837 =>  388,
      838 to   840 =>  389,
      841 to   842 =>  390,
      843 to   844 =>  391,
      845 to   847 =>  392,
      848 to   849 =>  393,
      850 to   852 =>  394,
      853 to   854 =>  395,
      855 to   856 =>  396,
      857 to   859 =>  397,
      860 to   861 =>  398,
      862 to   864 =>  399,
      865 to   866 =>  400,
      867 to   869 =>  401,
      870 to   871 =>  402,
      872 to   873 =>  403,
      874 to   876 =>  404,
      877 to   878 =>  405,
      879 to   881 =>  406,
      882 to   883 =>  407,
      884 to   885 =>  408,
      886 to   888 =>  409,
      889 to   890 =>  410,
      891 to   893 =>  411,
      894 to   895 =>  412,
      896 to   898 =>  413,
      899 to   900 =>  414,
      901 to   903 =>  415,
      904 to   905 =>  416,
      906 to   907 =>  417,
      908 to   910 =>  418,
      911 to   912 =>  419,
      913 to   915 =>  420,
      916 to   917 =>  421,
      918 to   920 =>  422,
      921 to   922 =>  423,
      923 to   925 =>  424,
      926 to   927 =>  425,
      928 to   930 =>  426,
      931 to   932 =>  427,
      933 to   935 =>  428,
      936 to   937 =>  429,
      938 to   939 =>  430,
      940 to   942 =>  431,
      943 to   944 =>  432,
      945 to   947 =>  433,
      948 to   949 =>  434,
      950 to   952 =>  435,
      953 to   954 =>  436,
      955 to   957 =>  437,
      958 to   959 =>  438,
      960 to   962 =>  439,
      963 to   964 =>  440,
      965 to   967 =>  441,
      968 to   969 =>  442,
      970 to   972 =>  443,
      973 to   974 =>  444,
      975 to   977 =>  445,
      978 to   979 =>  446,
      980 to   982 =>  447,
      983 to   985 =>  448,
      986 to   987 =>  449,
      988 to   990 =>  450,
      991 to   992 =>  451,
      993 to   995 =>  452,
      996 to   997 =>  453,
      998 to  1000 =>  454,
     1001 to  1002 =>  455,
     1003 to  1005 =>  456,
     1006 to  1007 =>  457,
     1008 to  1010 =>  458,
     1011 to  1012 =>  459,
     1013 to  1015 =>  460,
     1016 to  1018 =>  461,
     1019 to  1020 =>  462,
     1021 to  1023 =>  463,
     1024 to  1025 =>  464,
     1026 to  1028 =>  465,
     1029 to  1030 =>  466,
     1031 to  1033 =>  467,
     1034 to  1035 =>  468,
     1036 to  1038 =>  469,
     1039 to  1041 =>  470,
     1042 to  1043 =>  471,
     1044 to  1046 =>  472,
     1047 to  1048 =>  473,
     1049 to  1051 =>  474,
     1052 to  1054 =>  475,
     1055 to  1056 =>  476,
     1057 to  1059 =>  477,
     1060 to  1061 =>  478,
     1062 to  1064 =>  479,
     1065 to  1067 =>  480,
     1068 to  1069 =>  481,
     1070 to  1072 =>  482,
     1073 to  1074 =>  483,
     1075 to  1077 =>  484,
     1078 to  1080 =>  485,
     1081 to  1082 =>  486,
     1083 to  1085 =>  487,
     1086 to  1087 =>  488,
     1088 to  1090 =>  489,
     1091 to  1093 =>  490,
     1094 to  1095 =>  491,
     1096 to  1098 =>  492,
     1099 to  1101 =>  493,
     1102 to  1103 =>  494,
     1104 to  1106 =>  495,
     1107 to  1109 =>  496,
     1110 to  1111 =>  497,
     1112 to  1114 =>  498,
     1115 to  1116 =>  499,
     1117 to  1119 =>  500,
     1120 to  1122 =>  501,
     1123 to  1124 =>  502,
     1125 to  1127 =>  503,
     1128 to  1130 =>  504,
     1131 to  1132 =>  505,
     1133 to  1135 =>  506,
     1136 to  1138 =>  507,
     1139 to  1141 =>  508,
     1142 to  1143 =>  509,
     1144 to  1146 =>  510,
     1147 to  1149 =>  511,
     1150 to  1151 =>  512,
     1152 to  1154 =>  513,
     1155 to  1157 =>  514,
     1158 to  1159 =>  515,
     1160 to  1162 =>  516,
     1163 to  1165 =>  517,
     1166 to  1168 =>  518,
     1169 to  1170 =>  519,
     1171 to  1173 =>  520,
     1174 to  1176 =>  521,
     1177 to  1178 =>  522,
     1179 to  1181 =>  523,
     1182 to  1184 =>  524,
     1185 to  1187 =>  525,
     1188 to  1189 =>  526,
     1190 to  1192 =>  527,
     1193 to  1195 =>  528,
     1196 to  1198 =>  529,
     1199 to  1200 =>  530,
     1201 to  1203 =>  531,
     1204 to  1206 =>  532,
     1207 to  1209 =>  533,
     1210 to  1211 =>  534,
     1212 to  1214 =>  535,
     1215 to  1217 =>  536,
     1218 to  1220 =>  537,
     1221 to  1222 =>  538,
     1223 to  1225 =>  539,
     1226 to  1228 =>  540,
     1229 to  1231 =>  541,
     1232 to  1234 =>  542,
     1235 to  1236 =>  543,
     1237 to  1239 =>  544,
     1240 to  1242 =>  545,
     1243 to  1245 =>  546,
     1246 to  1248 =>  547,
     1249 to  1250 =>  548,
     1251 to  1253 =>  549,
     1254 to  1256 =>  550,
     1257 to  1259 =>  551,
     1260 to  1262 =>  552,
     1263 to  1265 =>  553,
     1266 to  1267 =>  554,
     1268 to  1270 =>  555,
     1271 to  1273 =>  556,
     1274 to  1276 =>  557,
     1277 to  1279 =>  558,
     1280 to  1282 =>  559,
     1283 to  1284 =>  560,
     1285 to  1287 =>  561,
     1288 to  1290 =>  562,
     1291 to  1293 =>  563,
     1294 to  1296 =>  564,
     1297 to  1299 =>  565,
     1300 to  1302 =>  566,
     1303 to  1304 =>  567,
     1305 to  1307 =>  568,
     1308 to  1310 =>  569,
     1311 to  1313 =>  570,
     1314 to  1316 =>  571,
     1317 to  1319 =>  572,
     1320 to  1322 =>  573,
     1323 to  1325 =>  574,
     1326 to  1328 =>  575,
     1329 to  1331 =>  576,
     1332 to  1333 =>  577,
     1334 to  1336 =>  578,
     1337 to  1339 =>  579,
     1340 to  1342 =>  580,
     1343 to  1345 =>  581,
     1346 to  1348 =>  582,
     1349 to  1351 =>  583,
     1352 to  1354 =>  584,
     1355 to  1357 =>  585,
     1358 to  1360 =>  586,
     1361 to  1363 =>  587,
     1364 to  1366 =>  588,
     1367 to  1369 =>  589,
     1370 to  1372 =>  590,
     1373 to  1375 =>  591,
     1376 to  1378 =>  592,
     1379 to  1381 =>  593,
     1382 to  1384 =>  594,
     1385 to  1387 =>  595,
     1388 to  1390 =>  596,
     1391 to  1393 =>  597,
     1394 to  1396 =>  598,
     1397 to  1399 =>  599,
     1400 to  1402 =>  600,
     1403 to  1405 =>  601,
     1406 to  1408 =>  602,
     1409 to  1411 =>  603,
     1412 to  1414 =>  604,
     1415 to  1417 =>  605,
     1418 to  1420 =>  606,
     1421 to  1423 =>  607,
     1424 to  1426 =>  608,
     1427 to  1429 =>  609,
     1430 to  1432 =>  610,
     1433 to  1435 =>  611,
     1436 to  1438 =>  612,
     1439 to  1441 =>  613,
     1442 to  1444 =>  614,
     1445 to  1447 =>  615,
     1448 to  1450 =>  616,
     1451 to  1453 =>  617,
     1454 to  1456 =>  618,
     1457 to  1460 =>  619,
     1461 to  1463 =>  620,
     1464 to  1466 =>  621,
     1467 to  1469 =>  622,
     1470 to  1472 =>  623,
     1473 to  1475 =>  624,
     1476 to  1478 =>  625,
     1479 to  1481 =>  626,
     1482 to  1484 =>  627,
     1485 to  1488 =>  628,
     1489 to  1491 =>  629,
     1492 to  1494 =>  630,
     1495 to  1497 =>  631,
     1498 to  1500 =>  632,
     1501 to  1503 =>  633,
     1504 to  1506 =>  634,
     1507 to  1510 =>  635,
     1511 to  1513 =>  636,
     1514 to  1516 =>  637,
     1517 to  1519 =>  638,
     1520 to  1522 =>  639,
     1523 to  1525 =>  640,
     1526 to  1529 =>  641,
     1530 to  1532 =>  642,
     1533 to  1535 =>  643,
     1536 to  1538 =>  644,
     1539 to  1541 =>  645,
     1542 to  1545 =>  646,
     1546 to  1548 =>  647,
     1549 to  1551 =>  648,
     1552 to  1554 =>  649,
     1555 to  1558 =>  650,
     1559 to  1561 =>  651,
     1562 to  1564 =>  652,
     1565 to  1567 =>  653,
     1568 to  1570 =>  654,
     1571 to  1574 =>  655,
     1575 to  1577 =>  656,
     1578 to  1580 =>  657,
     1581 to  1584 =>  658,
     1585 to  1587 =>  659,
     1588 to  1590 =>  660,
     1591 to  1593 =>  661,
     1594 to  1597 =>  662,
     1598 to  1600 =>  663,
     1601 to  1603 =>  664,
     1604 to  1607 =>  665,
     1608 to  1610 =>  666,
     1611 to  1613 =>  667,
     1614 to  1617 =>  668,
     1618 to  1620 =>  669,
     1621 to  1623 =>  670,
     1624 to  1627 =>  671,
     1628 to  1630 =>  672,
     1631 to  1633 =>  673,
     1634 to  1637 =>  674,
     1638 to  1640 =>  675,
     1641 to  1643 =>  676,
     1644 to  1647 =>  677,
     1648 to  1650 =>  678,
     1651 to  1653 =>  679,
     1654 to  1657 =>  680,
     1658 to  1660 =>  681,
     1661 to  1664 =>  682,
     1665 to  1667 =>  683,
     1668 to  1670 =>  684,
     1671 to  1674 =>  685,
     1675 to  1677 =>  686,
     1678 to  1681 =>  687,
     1682 to  1684 =>  688,
     1685 to  1688 =>  689,
     1689 to  1691 =>  690,
     1692 to  1694 =>  691,
     1695 to  1698 =>  692,
     1699 to  1701 =>  693,
     1702 to  1705 =>  694,
     1706 to  1708 =>  695,
     1709 to  1712 =>  696,
     1713 to  1715 =>  697,
     1716 to  1719 =>  698,
     1720 to  1722 =>  699,
     1723 to  1726 =>  700,
     1727 to  1729 =>  701,
     1730 to  1733 =>  702,
     1734 to  1736 =>  703,
     1737 to  1740 =>  704,
     1741 to  1743 =>  705,
     1744 to  1747 =>  706,
     1748 to  1750 =>  707,
     1751 to  1754 =>  708,
     1755 to  1758 =>  709,
     1759 to  1761 =>  710,
     1762 to  1765 =>  711,
     1766 to  1768 =>  712,
     1769 to  1772 =>  713,
     1773 to  1775 =>  714,
     1776 to  1779 =>  715,
     1780 to  1783 =>  716,
     1784 to  1786 =>  717,
     1787 to  1790 =>  718,
     1791 to  1793 =>  719,
     1794 to  1797 =>  720,
     1798 to  1801 =>  721,
     1802 to  1804 =>  722,
     1805 to  1808 =>  723,
     1809 to  1812 =>  724,
     1813 to  1815 =>  725,
     1816 to  1819 =>  726,
     1820 to  1823 =>  727,
     1824 to  1826 =>  728,
     1827 to  1830 =>  729,
     1831 to  1834 =>  730,
     1835 to  1837 =>  731,
     1838 to  1841 =>  732,
     1842 to  1845 =>  733,
     1846 to  1848 =>  734,
     1849 to  1852 =>  735,
     1853 to  1856 =>  736,
     1857 to  1860 =>  737,
     1861 to  1863 =>  738,
     1864 to  1867 =>  739,
     1868 to  1871 =>  740,
     1872 to  1875 =>  741,
     1876 to  1878 =>  742,
     1879 to  1882 =>  743,
     1883 to  1886 =>  744,
     1887 to  1890 =>  745,
     1891 to  1894 =>  746,
     1895 to  1897 =>  747,
     1898 to  1901 =>  748,
     1902 to  1905 =>  749,
     1906 to  1909 =>  750,
     1910 to  1913 =>  751,
     1914 to  1916 =>  752,
     1917 to  1920 =>  753,
     1921 to  1924 =>  754,
     1925 to  1928 =>  755,
     1929 to  1932 =>  756,
     1933 to  1936 =>  757,
     1937 to  1940 =>  758,
     1941 to  1944 =>  759,
     1945 to  1947 =>  760,
     1948 to  1951 =>  761,
     1952 to  1955 =>  762,
     1956 to  1959 =>  763,
     1960 to  1963 =>  764,
     1964 to  1967 =>  765,
     1968 to  1971 =>  766,
     1972 to  1975 =>  767,
     1976 to  1979 =>  768,
     1980 to  1983 =>  769,
     1984 to  1987 =>  770,
     1988 to  1991 =>  771,
     1992 to  1995 =>  772,
     1996 to  1999 =>  773,
     2000 to  2003 =>  774,
     2004 to  2007 =>  775,
     2008 to  2011 =>  776,
     2012 to  2015 =>  777,
     2016 to  2019 =>  778,
     2020 to  2023 =>  779,
     2024 to  2027 =>  780,
     2028 to  2031 =>  781,
     2032 to  2035 =>  782,
     2036 to  2039 =>  783,
     2040 to  2043 =>  784,
     2044 to  2047 =>  785,
     2048 to  2052 =>  786,
     2053 to  2056 =>  787,
     2057 to  2060 =>  788,
     2061 to  2064 =>  789,
     2065 to  2068 =>  790,
     2069 to  2072 =>  791,
     2073 to  2076 =>  792,
     2077 to  2080 =>  793,
     2081 to  2085 =>  794,
     2086 to  2089 =>  795,
     2090 to  2093 =>  796,
     2094 to  2097 =>  797,
     2098 to  2101 =>  798,
     2102 to  2106 =>  799,
     2107 to  2110 =>  800,
     2111 to  2114 =>  801,
     2115 to  2118 =>  802,
     2119 to  2123 =>  803,
     2124 to  2127 =>  804,
     2128 to  2131 =>  805,
     2132 to  2135 =>  806,
     2136 to  2140 =>  807,
     2141 to  2144 =>  808,
     2145 to  2148 =>  809,
     2149 to  2152 =>  810,
     2153 to  2157 =>  811,
     2158 to  2161 =>  812,
     2162 to  2165 =>  813,
     2166 to  2170 =>  814,
     2171 to  2174 =>  815,
     2175 to  2179 =>  816,
     2180 to  2183 =>  817,
     2184 to  2187 =>  818,
     2188 to  2192 =>  819,
     2193 to  2196 =>  820,
     2197 to  2200 =>  821,
     2201 to  2205 =>  822,
     2206 to  2209 =>  823,
     2210 to  2214 =>  824,
     2215 to  2218 =>  825,
     2219 to  2223 =>  826,
     2224 to  2227 =>  827,
     2228 to  2232 =>  828,
     2233 to  2236 =>  829,
     2237 to  2241 =>  830,
     2242 to  2245 =>  831,
     2246 to  2250 =>  832,
     2251 to  2254 =>  833,
     2255 to  2259 =>  834,
     2260 to  2263 =>  835,
     2264 to  2268 =>  836,
     2269 to  2272 =>  837,
     2273 to  2277 =>  838,
     2278 to  2282 =>  839,
     2283 to  2286 =>  840,
     2287 to  2291 =>  841,
     2292 to  2295 =>  842,
     2296 to  2300 =>  843,
     2301 to  2305 =>  844,
     2306 to  2309 =>  845,
     2310 to  2314 =>  846,
     2315 to  2319 =>  847,
     2320 to  2323 =>  848,
     2324 to  2328 =>  849,
     2329 to  2333 =>  850,
     2334 to  2337 =>  851,
     2338 to  2342 =>  852,
     2343 to  2347 =>  853,
     2348 to  2352 =>  854,
     2353 to  2356 =>  855,
     2357 to  2361 =>  856,
     2362 to  2366 =>  857,
     2367 to  2371 =>  858,
     2372 to  2375 =>  859,
     2376 to  2380 =>  860,
     2381 to  2385 =>  861,
     2386 to  2390 =>  862,
     2391 to  2395 =>  863,
     2396 to  2400 =>  864,
     2401 to  2404 =>  865,
     2405 to  2409 =>  866,
     2410 to  2414 =>  867,
     2415 to  2419 =>  868,
     2420 to  2424 =>  869,
     2425 to  2429 =>  870,
     2430 to  2434 =>  871,
     2435 to  2439 =>  872,
     2440 to  2444 =>  873,
     2445 to  2449 =>  874,
     2450 to  2454 =>  875,
     2455 to  2459 =>  876,
     2460 to  2464 =>  877,
     2465 to  2469 =>  878,
     2470 to  2474 =>  879,
     2475 to  2479 =>  880,
     2480 to  2484 =>  881,
     2485 to  2489 =>  882,
     2490 to  2494 =>  883,
     2495 to  2499 =>  884,
     2500 to  2504 =>  885,
     2505 to  2509 =>  886,
     2510 to  2515 =>  887,
     2516 to  2520 =>  888,
     2521 to  2525 =>  889,
     2526 to  2530 =>  890,
     2531 to  2535 =>  891,
     2536 to  2540 =>  892,
     2541 to  2546 =>  893,
     2547 to  2551 =>  894,
     2552 to  2556 =>  895,
     2557 to  2561 =>  896,
     2562 to  2567 =>  897,
     2568 to  2572 =>  898,
     2573 to  2577 =>  899,
     2578 to  2582 =>  900,
     2583 to  2588 =>  901,
     2589 to  2593 =>  902,
     2594 to  2598 =>  903,
     2599 to  2604 =>  904,
     2605 to  2609 =>  905,
     2610 to  2615 =>  906,
     2616 to  2620 =>  907,
     2621 to  2625 =>  908,
     2626 to  2631 =>  909,
     2632 to  2636 =>  910,
     2637 to  2642 =>  911,
     2643 to  2647 =>  912,
     2648 to  2653 =>  913,
     2654 to  2658 =>  914,
     2659 to  2664 =>  915,
     2665 to  2669 =>  916,
     2670 to  2675 =>  917,
     2676 to  2680 =>  918,
     2681 to  2686 =>  919,
     2687 to  2691 =>  920,
     2692 to  2697 =>  921,
     2698 to  2703 =>  922,
     2704 to  2708 =>  923,
     2709 to  2714 =>  924,
     2715 to  2719 =>  925,
     2720 to  2725 =>  926,
     2726 to  2731 =>  927,
     2732 to  2737 =>  928,
     2738 to  2742 =>  929,
     2743 to  2748 =>  930,
     2749 to  2754 =>  931,
     2755 to  2759 =>  932,
     2760 to  2765 =>  933,
     2766 to  2771 =>  934,
     2772 to  2777 =>  935,
     2778 to  2783 =>  936,
     2784 to  2789 =>  937,
     2790 to  2794 =>  938,
     2795 to  2800 =>  939,
     2801 to  2806 =>  940,
     2807 to  2812 =>  941,
     2813 to  2818 =>  942,
     2819 to  2824 =>  943,
     2825 to  2830 =>  944,
     2831 to  2836 =>  945,
     2837 to  2842 =>  946,
     2843 to  2848 =>  947,
     2849 to  2854 =>  948,
     2855 to  2860 =>  949,
     2861 to  2866 =>  950,
     2867 to  2872 =>  951,
     2873 to  2878 =>  952,
     2879 to  2884 =>  953,
     2885 to  2890 =>  954,
     2891 to  2896 =>  955,
     2897 to  2903 =>  956,
     2904 to  2909 =>  957,
     2910 to  2915 =>  958,
     2916 to  2921 =>  959,
     2922 to  2927 =>  960,
     2928 to  2934 =>  961,
     2935 to  2940 =>  962,
     2941 to  2946 =>  963,
     2947 to  2952 =>  964,
     2953 to  2959 =>  965,
     2960 to  2965 =>  966,
     2966 to  2971 =>  967,
     2972 to  2978 =>  968,
     2979 to  2984 =>  969,
     2985 to  2991 =>  970,
     2992 to  2997 =>  971,
     2998 to  3004 =>  972,
     3005 to  3010 =>  973,
     3011 to  3016 =>  974,
     3017 to  3023 =>  975,
     3024 to  3030 =>  976,
     3031 to  3036 =>  977,
     3037 to  3043 =>  978,
     3044 to  3049 =>  979,
     3050 to  3056 =>  980,
     3057 to  3062 =>  981,
     3063 to  3069 =>  982,
     3070 to  3076 =>  983,
     3077 to  3082 =>  984,
     3083 to  3089 =>  985,
     3090 to  3096 =>  986,
     3097 to  3103 =>  987,
     3104 to  3109 =>  988,
     3110 to  3116 =>  989,
     3117 to  3123 =>  990,
     3124 to  3130 =>  991,
     3131 to  3137 =>  992,
     3138 to  3143 =>  993,
     3144 to  3150 =>  994,
     3151 to  3157 =>  995,
     3158 to  3164 =>  996,
     3165 to  3171 =>  997,
     3172 to  3178 =>  998,
     3179 to  3185 =>  999,
     3186 to  3192 => 1000,
     3193 to  3199 => 1001,
     3200 to  3206 => 1002,
     3207 to  3213 => 1003,
     3214 to  3220 => 1004,
     3221 to  3227 => 1005,
     3228 to  3235 => 1006,
     3236 to  3242 => 1007,
     3243 to  3249 => 1008,
     3250 to  3256 => 1009,
     3257 to  3263 => 1010,
     3264 to  3271 => 1011,
     3272 to  3278 => 1012,
     3279 to  3285 => 1013,
     3286 to  3293 => 1014,
     3294 to  3300 => 1015,
     3301 to  3307 => 1016,
     3308 to  3315 => 1017,
     3316 to  3322 => 1018,
     3323 to  3330 => 1019,
     3331 to  3337 => 1020,
     3338 to  3345 => 1021,
     3346 to  3352 => 1022,
     3353 to  3360 => 1023,
     3361 to  3367 => 1024,
     3368 to  3375 => 1025,
     3376 to  3383 => 1026,
     3384 to  3390 => 1027,
     3391 to  3398 => 1028,
     3399 to  3406 => 1029,
     3407 to  3413 => 1030,
     3414 to  3421 => 1031,
     3422 to  3429 => 1032,
     3430 to  3437 => 1033,
     3438 to  3444 => 1034,
     3445 to  3452 => 1035,
     3453 to  3460 => 1036,
     3461 to  3468 => 1037,
     3469 to  3476 => 1038,
     3477 to  3484 => 1039,
     3485 to  3492 => 1040,
     3493 to  3500 => 1041,
     3501 to  3508 => 1042,
     3509 to  3516 => 1043,
     3517 to  3524 => 1044,
     3525 to  3532 => 1045,
     3533 to  3541 => 1046,
     3542 to  3549 => 1047,
     3550 to  3557 => 1048,
     3558 to  3565 => 1049,
     3566 to  3573 => 1050,
     3574 to  3582 => 1051,
     3583 to  3590 => 1052,
     3591 to  3598 => 1053,
     3599 to  3607 => 1054,
     3608 to  3615 => 1055,
     3616 to  3624 => 1056,
     3625 to  3632 => 1057,
     3633 to  3641 => 1058,
     3642 to  3649 => 1059,
     3650 to  3658 => 1060,
     3659 to  3666 => 1061,
     3667 to  3675 => 1062,
     3676 to  3684 => 1063,
     3685 to  3692 => 1064,
     3693 to  3701 => 1065,
     3702 to  3710 => 1066,
     3711 to  3719 => 1067,
     3720 to  3727 => 1068,
     3728 to  3736 => 1069,
     3737 to  3745 => 1070,
     3746 to  3754 => 1071,
     3755 to  3763 => 1072,
     3764 to  3772 => 1073,
     3773 to  3781 => 1074,
     3782 to  3790 => 1075,
     3791 to  3799 => 1076,
     3800 to  3808 => 1077,
     3809 to  3817 => 1078,
     3818 to  3827 => 1079,
     3828 to  3836 => 1080,
     3837 to  3845 => 1081,
     3846 to  3854 => 1082,
     3855 to  3864 => 1083,
     3865 to  3873 => 1084,
     3874 to  3882 => 1085,
     3883 to  3892 => 1086,
     3893 to  3901 => 1087,
     3902 to  3911 => 1088,
     3912 to  3920 => 1089,
     3921 to  3930 => 1090,
     3931 to  3940 => 1091,
     3941 to  3949 => 1092,
     3950 to  3959 => 1093,
     3960 to  3969 => 1094,
     3970 to  3978 => 1095,
     3979 to  3988 => 1096,
     3989 to  3998 => 1097,
     3999 to  4008 => 1098,
     4009 to  4018 => 1099,
     4019 to  4028 => 1100,
     4029 to  4038 => 1101,
     4039 to  4048 => 1102,
     4049 to  4058 => 1103,
     4059 to  4068 => 1104,
     4069 to  4078 => 1105,
     4079 to  4088 => 1106,
     4089 to  4099 => 1107,
     4100 to  4109 => 1108,
     4110 to  4119 => 1109,
     4120 to  4130 => 1110,
     4131 to  4140 => 1111,
     4141 to  4150 => 1112,
     4151 to  4161 => 1113,
     4162 to  4171 => 1114,
     4172 to  4182 => 1115,
     4183 to  4193 => 1116,
     4194 to  4203 => 1117,
     4204 to  4214 => 1118,
     4215 to  4225 => 1119,
     4226 to  4235 => 1120,
     4236 to  4246 => 1121,
     4247 to  4257 => 1122,
     4258 to  4268 => 1123,
     4269 to  4279 => 1124,
     4280 to  4290 => 1125,
     4291 to  4301 => 1126,
     4302 to  4312 => 1127,
     4313 to  4323 => 1128,
     4324 to  4335 => 1129,
     4336 to  4346 => 1130,
     4347 to  4357 => 1131,
     4358 to  4369 => 1132,
     4370 to  4380 => 1133,
     4381 to  4391 => 1134,
     4392 to  4403 => 1135,
     4404 to  4414 => 1136,
     4415 to  4426 => 1137,
     4427 to  4438 => 1138,
     4439 to  4449 => 1139,
     4450 to  4461 => 1140,
     4462 to  4473 => 1141,
     4474 to  4485 => 1142,
     4486 to  4497 => 1143,
     4498 to  4509 => 1144,
     4510 to  4521 => 1145,
     4522 to  4533 => 1146,
     4534 to  4545 => 1147,
     4546 to  4557 => 1148,
     4558 to  4569 => 1149,
     4570 to  4581 => 1150,
     4582 to  4594 => 1151,
     4595 to  4606 => 1152,
     4607 to  4619 => 1153,
     4620 to  4631 => 1154,
     4632 to  4644 => 1155,
     4645 to  4656 => 1156,
     4657 to  4669 => 1157,
     4670 to  4682 => 1158,
     4683 to  4694 => 1159,
     4695 to  4707 => 1160,
     4708 to  4720 => 1161,
     4721 to  4733 => 1162,
     4734 to  4746 => 1163,
     4747 to  4759 => 1164,
     4760 to  4772 => 1165,
     4773 to  4786 => 1166,
     4787 to  4799 => 1167,
     4800 to  4812 => 1168,
     4813 to  4826 => 1169,
     4827 to  4839 => 1170,
     4840 to  4853 => 1171,
     4854 to  4866 => 1172,
     4867 to  4880 => 1173,
     4881 to  4893 => 1174,
     4894 to  4907 => 1175,
     4908 to  4921 => 1176,
     4922 to  4935 => 1177,
     4936 to  4949 => 1178,
     4950 to  4963 => 1179,
     4964 to  4977 => 1180,
     4978 to  4991 => 1181,
     4992 to  5006 => 1182,
     5007 to  5020 => 1183,
     5021 to  5034 => 1184,
     5035 to  5049 => 1185,
     5050 to  5063 => 1186,
     5064 to  5078 => 1187,
     5079 to  5093 => 1188,
     5094 to  5107 => 1189,
     5108 to  5122 => 1190,
     5123 to  5137 => 1191,
     5138 to  5152 => 1192,
     5153 to  5167 => 1193,
     5168 to  5182 => 1194,
     5183 to  5197 => 1195,
     5198 to  5213 => 1196,
     5214 to  5228 => 1197,
     5229 to  5243 => 1198,
     5244 to  5259 => 1199,
     5260 to  5275 => 1200,
     5276 to  5290 => 1201,
     5291 to  5306 => 1202,
     5307 to  5322 => 1203,
     5323 to  5338 => 1204,
     5339 to  5354 => 1205,
     5355 to  5370 => 1206,
     5371 to  5386 => 1207,
     5387 to  5402 => 1208,
     5403 to  5419 => 1209,
     5420 to  5435 => 1210,
     5436 to  5452 => 1211,
     5453 to  5468 => 1212,
     5469 to  5485 => 1213,
     5486 to  5502 => 1214,
     5503 to  5519 => 1215,
     5520 to  5536 => 1216,
     5537 to  5553 => 1217,
     5554 to  5570 => 1218,
     5571 to  5587 => 1219,
     5588 to  5604 => 1220,
     5605 to  5622 => 1221,
     5623 to  5639 => 1222,
     5640 to  5657 => 1223,
     5658 to  5675 => 1224,
     5676 to  5693 => 1225,
     5694 to  5710 => 1226,
     5711 to  5728 => 1227,
     5729 to  5747 => 1228,
     5748 to  5765 => 1229,
     5766 to  5783 => 1230,
     5784 to  5802 => 1231,
     5803 to  5820 => 1232,
     5821 to  5839 => 1233,
     5840 to  5858 => 1234,
     5859 to  5876 => 1235,
     5877 to  5895 => 1236,
     5896 to  5914 => 1237,
     5915 to  5934 => 1238,
     5935 to  5953 => 1239,
     5954 to  5972 => 1240,
     5973 to  5992 => 1241,
     5993 to  6012 => 1242,
     6013 to  6031 => 1243,
     6032 to  6051 => 1244,
     6052 to  6071 => 1245,
     6072 to  6091 => 1246,
     6092 to  6112 => 1247,
     6113 to  6132 => 1248,
     6133 to  6152 => 1249,
     6153 to  6173 => 1250,
     6174 to  6194 => 1251,
     6195 to  6214 => 1252,
     6215 to  6235 => 1253,
     6236 to  6257 => 1254,
     6258 to  6278 => 1255,
     6279 to  6299 => 1256,
     6300 to  6321 => 1257,
     6322 to  6342 => 1258,
     6343 to  6364 => 1259,
     6365 to  6386 => 1260,
     6387 to  6408 => 1261,
     6409 to  6430 => 1262,
     6431 to  6452 => 1263,
     6453 to  6475 => 1264,
     6476 to  6498 => 1265,
     6499 to  6520 => 1266,
     6521 to  6543 => 1267,
     6544 to  6566 => 1268,
     6567 to  6589 => 1269,
     6590 to  6613 => 1270,
     6614 to  6636 => 1271,
     6637 to  6660 => 1272,
     6661 to  6684 => 1273,
     6685 to  6708 => 1274,
     6709 to  6732 => 1275,
     6733 to  6756 => 1276,
     6757 to  6780 => 1277,
     6781 to  6805 => 1278,
     6806 to  6830 => 1279,
     6831 to  6855 => 1280,
     6856 to  6880 => 1281,
     6881 to  6905 => 1282,
     6906 to  6930 => 1283,
     6931 to  6956 => 1284,
     6957 to  6982 => 1285,
     6983 to  7008 => 1286,
     7009 to  7034 => 1287,
     7035 to  7060 => 1288,
     7061 to  7087 => 1289,
     7088 to  7113 => 1290,
     7114 to  7140 => 1291,
     7141 to  7167 => 1292,
     7168 to  7194 => 1293,
     7195 to  7222 => 1294,
     7223 to  7249 => 1295,
     7250 to  7277 => 1296,
     7278 to  7305 => 1297,
     7306 to  7333 => 1298,
     7334 to  7362 => 1299,
     7363 to  7390 => 1300,
     7391 to  7419 => 1301,
     7420 to  7448 => 1302,
     7449 to  7478 => 1303,
     7479 to  7507 => 1304,
     7508 to  7537 => 1305,
     7538 to  7567 => 1306,
     7568 to  7597 => 1307,
     7598 to  7627 => 1308,
     7628 to  7658 => 1309,
     7659 to  7688 => 1310,
     7689 to  7720 => 1311,
     7721 to  7751 => 1312,
     7752 to  7782 => 1313,
     7783 to  7814 => 1314,
     7815 to  7846 => 1315,
     7847 to  7878 => 1316,
     7879 to  7911 => 1317,
     7912 to  7944 => 1318,
     7945 to  7976 => 1319,
     7977 to  8010 => 1320,
     8011 to  8043 => 1321,
     8044 to  8077 => 1322,
     8078 to  8111 => 1323,
     8112 to  8145 => 1324,
     8146 to  8180 => 1325,
     8181 to  8215 => 1326,
     8216 to  8250 => 1327,
     8251 to  8285 => 1328,
     8286 to  8321 => 1329,
     8322 to  8357 => 1330,
     8358 to  8393 => 1331,
     8394 to  8430 => 1332,
     8431 to  8467 => 1333,
     8468 to  8504 => 1334,
     8505 to  8542 => 1335,
     8543 to  8580 => 1336,
     8581 to  8618 => 1337,
     8619 to  8656 => 1338,
     8657 to  8695 => 1339,
     8696 to  8734 => 1340,
     8735 to  8774 => 1341,
     8775 to  8813 => 1342,
     8814 to  8854 => 1343,
     8855 to  8894 => 1344,
     8895 to  8935 => 1345,
     8936 to  8976 => 1346,
     8977 to  9018 => 1347,
     9019 to  9060 => 1348,
     9061 to  9102 => 1349,
     9103 to  9145 => 1350,
     9146 to  9188 => 1351,
     9189 to  9231 => 1352,
     9232 to  9275 => 1353,
     9276 to  9319 => 1354,
     9320 to  9364 => 1355,
     9365 to  9409 => 1356,
     9410 to  9455 => 1357,
     9456 to  9501 => 1358,
     9502 to  9547 => 1359,
     9548 to  9594 => 1360,
     9595 to  9641 => 1361,
     9642 to  9689 => 1362,
     9690 to  9737 => 1363,
     9738 to  9785 => 1364,
     9786 to  9834 => 1365,
     9835 to  9884 => 1366,
     9885 to  9934 => 1367,
     9935 to  9984 => 1368,
     9985 to 10035 => 1369,
    10036 to 10087 => 1370,
    10088 to 10139 => 1371,
    10140 to 10191 => 1372,
    10192 to 10244 => 1373,
    10245 to 10298 => 1374,
    10299 to 10352 => 1375,
    10353 to 10407 => 1376,
    10408 to 10462 => 1377,
    10463 to 10518 => 1378,
    10519 to 10574 => 1379,
    10575 to 10631 => 1380,
    10632 to 10689 => 1381,
    10690 to 10747 => 1382,
    10748 to 10805 => 1383,
    10806 to 10865 => 1384,
    10866 to 10925 => 1385,
    10926 to 10986 => 1386,
    10987 to 11047 => 1387,
    11048 to 11109 => 1388,
    11110 to 11171 => 1389,
    11172 to 11235 => 1390,
    11236 to 11299 => 1391,
    11300 to 11364 => 1392,
    11365 to 11429 => 1393,
    11430 to 11495 => 1394,
    11496 to 11562 => 1395,
    11563 to 11630 => 1396,
    11631 to 11698 => 1397,
    11699 to 11768 => 1398,
    11769 to 11838 => 1399,
    11839 to 11909 => 1400,
    11910 to 11980 => 1401,
    11981 to 12053 => 1402,
    12054 to 12126 => 1403,
    12127 to 12201 => 1404,
    12202 to 12276 => 1405,
    12277 to 12352 => 1406,
    12353 to 12429 => 1407,
    12430 to 12507 => 1408,
    12508 to 12586 => 1409,
    12587 to 12666 => 1410,
    12667 to 12747 => 1411,
    12748 to 12829 => 1412,
    12830 to 12912 => 1413,
    12913 to 12996 => 1414,
    12997 to 13081 => 1415,
    13082 to 13167 => 1416,
    13168 to 13254 => 1417,
    13255 to 13342 => 1418,
    13343 to 13432 => 1419,
    13433 to 13523 => 1420,
    13524 to 13615 => 1421,
    13616 to 13708 => 1422,
    13709 to 13802 => 1423,
    13803 to 13898 => 1424,
    13899 to 13995 => 1425,
    13996 to 14094 => 1426,
    14095 to 14193 => 1427,
    14194 to 14294 => 1428,
    14295 to 14397 => 1429,
    14398 to 14501 => 1430,
    14502 to 14606 => 1431,
    14607 to 14713 => 1432,
    14714 to 14822 => 1433,
    14823 to 14932 => 1434,
    14933 to 15044 => 1435,
    15045 to 15157 => 1436,
    15158 to 15272 => 1437,
    15273 to 15389 => 1438,
    15390 to 15508 => 1439,
    15509 to 15628 => 1440,
    15629 to 15750 => 1441,
    15751 to 15875 => 1442,
    15876 to 16001 => 1443,
    16002 to 16129 => 1444,
    16130 to 16259 => 1445,
    16260 to 16391 => 1446,
    16392 to 16525 => 1447,
    16526 to 16662 => 1448,
    16663 to 16801 => 1449,
    16802 to 16942 => 1450,
    16943 to 17085 => 1451,
    17086 to 17231 => 1452,
    17232 to 17379 => 1453,
    17380 to 17530 => 1454,
    17531 to 17683 => 1455,
    17684 to 17840 => 1456,
    17841 to 17998 => 1457,
    17999 to 18160 => 1458,
    18161 to 18325 => 1459,
    18326 to 18492 => 1460,
    18493 to 18663 => 1461,
    18664 to 18836 => 1462,
    18837 to 19013 => 1463,
    19014 to 19194 => 1464,
    19195 to 19377 => 1465,
    19378 to 19565 => 1466,
    19566 to 19755 => 1467,
    19756 to 19950 => 1468,
    19951 to 20148 => 1469,
    20149 to 20350 => 1470,
    20351 to 20557 => 1471,
    20558 to 20767 => 1472,
    20768 to 20982 => 1473,
    20983 to 21201 => 1474,
    21202 to 21425 => 1475,
    21426 to 21654 => 1476,
    21655 to 21887 => 1477,
    21888 to 22126 => 1478,
    22127 to 22370 => 1479,
    22371 to 22619 => 1480,
    22620 to 22874 => 1481,
    22875 to 23134 => 1482,
    23135 to 23400 => 1483,
    23401 to 23673 => 1484,
    23674 to 23952 => 1485,
    23953 to 24238 => 1486,
    24239 to 24530 => 1487,
    24531 to 24829 => 1488,
    24830 to 25136 => 1489,
    25137 to 25451 => 1490,
    25452 to 25773 => 1491,
    25774 to 26104 => 1492,
    26105 to 26443 => 1493,
    26444 to 26791 => 1494,
    26792 to 27148 => 1495,
    27149 to 27515 => 1496,
    27516 to 27892 => 1497,
    27893 to 28279 => 1498,
    28280 to 28677 => 1499,
    28678 to 29086 => 1500,
    29087 to 29507 => 1501,
    29508 to 29941 => 1502,
    29942 to 30387 => 1503,
    30388 to 30847 => 1504,
    30848 to 31321 => 1505,
    31322 to 31810 => 1506,
    31811 to 32314 => 1507,
    32315 to 32834 => 1508,
    32835 to 33371 => 1509,
    33372 to 33926 => 1510,
    33927 to 34499 => 1511,
    34500 to 35093 => 1512,
    35094 to 35707 => 1513,
    35708 to 36342 => 1514,
    36343 to 37001 => 1515,
    37002 to 37684 => 1516,
    37685 to 38393 => 1517,
    38394 to 39128 => 1518,
    39129 to 39893 => 1519,
    39894 to 40687 => 1520,
    40688 to 41514 => 1521,
    41515 to 42375 => 1522,
    42376 to 43273 => 1523,
    43274 to 44209 => 1524,
    44210 to 45187 => 1525,
    45188 to 46209 => 1526,
    46210 to 47278 => 1527,
    47279 to 48397 => 1528,
    48398 to 49571 => 1529,
    49572 to 50803 => 1530,
    50804 to 52097 => 1531,
    52098 to 53460 => 1532,
    53461 to 54895 => 1533,
    54896 to 56409 => 1534,
    56410 to 58010 => 1535,
    58011 to 59703 => 1536,
    59704 to 61498 => 1537,
    61499 to 63405 => 1538,
    63406 to 65433 => 1539,
    65434 to 67596 => 1540,
    67597 to 69906 => 1541,
    69907 to 72379 => 1542,
    72380 to 75034 => 1543,
    75035 to 77891 => 1544,
    77892 to 80974 => 1545,
    80975 to 84311 => 1546,
    84312 to 87934 => 1547,
    87935 to 91884 => 1548,
    91885 to 96204 => 1549,
    96205 to 100951 => 1550,
    100952 to 106191 => 1551,
    106192 to 112005 => 1552,
    112006 to 118493 => 1553,
    118494 to 125779 => 1554,
    125780 to 134020 => 1555,
    134021 to 143418 => 1556,
    143419 to 154236 => 1557,
    154237 to 166820 => 1558,
    166821 to 181645 => 1559,
    181646 to 199368 => 1560,
    199369 to 220934 => 1561,
    220935 to 247749 => 1562,
    247750 to 282008 => 1563,
    282009 to 327328 => 1564,
    327329 to 390156 => 1565,
    390157 to 483227 => 1566,
    483228 to 635926 => 1567,
    635927 to 732387 => 1568
  );

 end package roi_atan;
