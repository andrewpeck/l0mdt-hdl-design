//--------------------------------------------------------------------------------
//--  Department of Physics and Astronomy, UCI
//--  Priya Sundararajan
//--  priya.sundararajan@cern.ch
//--------------------------------------------------------------------------------
//--  Project: ATLAS L0MDT Trigger
//--  Description:
//--
//--------------------------------------------------------------------------------
//--  Revisions:
//--
//--------------------------------------------------------------------------------


////////////////////////////////////////////////////////////////////////////////////////////////////
// autogenerated file
// created by tb create on: 03-Jun-2020 (10:30:39)
// created by tb create for test: mtc
////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
`default_nettype wire
//`include "l0mdt_buses_constants.svh"

  module TopLevel_mtc #(
			parameter SLCPIPELINE_WIDTH = PL2MTC_LEN,
			parameter PTCALC_LEN = PTCALC2MTC_LEN,
			parameter MTC_LEN = MTC2SL_LEN,
			parameter TOTAL_PTCALC_BLKS=3,
			parameter MAX_MTC_PER_BCID=3,
    parameter DATA_WIDTH = 81,
    parameter FIFO_DEPTH = 6,
    parameter N_OUTPUTS = 3,
    parameter N_INPUTS = 3

) (
    input wire 			       clock,
    input wire 			       reset_n,
    input wire [SLCPIPELINE_WIDTH-1:0] slcpipeline [MAX_MTC_PER_BCID],
   // input wire 			       slcpipeline_vld [MAX_MTC_PER_BCID],
    input wire [PTCALC_LEN-1:0] 	       ptcalc [TOTAL_PTCALC_BLKS],
    input wire [1:0] 		       ptcalc_sel[TOTAL_PTCALC_BLKS],
    output wire [MTC_LEN-1:0] 	       mtc [MAX_MTC_PER_BCID],
    output wire 		       mtc_valid [MAX_MTC_PER_BCID]
);
   wire [MTC_LEN-1:0] 		       mtc_out [MAX_MTC_PER_BCID];
   wire 			       mtc_out_valid [MAX_MTC_PER_BCID];
   genvar 			       i;
   //Having issues monitoring buses >192 bits



     for( i=0; i<TOTAL_PTCALC_BLKS;i++)
       begin
	  assign ptcalc_sel[i] = i;

       end

   for( i=0; i<MAX_MTC_PER_BCID;i++)
       begin
	  assign slcpipeline[i]        = 0;
	  assign mtc_valid[i]          = mtc_out[i][MTC_LEN-1];

       end


   always@(posedge clock)
     begin
//	if(mtc_out[0][MTC_LEN-1] == 1)
//	  $display("TESTBENCH VAL MTC_OUT = 0x%x",mtc_out[0]);

     end

    //
    // Here define the signals to connect the input and output Spy+FIFO
    // blocks with the input and output of the DUT.
    // Here we define one for each of the FIFO signals, but the test
    // creator should remove unnecessary signals.
    //




    //
    // Here place the DUT block(s)
    //

    //Verilog Model
   mtc_builder_verilog#(
		   .PTCALC_WIDTH(PTCALC_LEN),
		    .SLCPIPELINE_WIDTH(SLCPIPELINE_WIDTH),
		    .TOTAL_PTCALC_BLKS(TOTAL_PTCALC_BLKS),
        .n_PRIMARY_MTC(3)
		    )
   mtc_builder_inst(
    		    .clock(clock),
		    .rst(~reset_n),
		    .srst(~reset_n),
		    .ptcalc(ptcalc),
		  //  .ptcalc_sel(ptcalc_sel),
		    .slcpipeline(slcpipeline),
		  //  .slcpipeline_vld(slcpipeline_vld),
		    .mtc(mtc_out)
		    //.mtc_valid(mtc_out_valid)
//    output logic [MTC_WIDTH:0] 	      mtc
    );


/*
   //VHDL Wrapper
   mtc_builder mtc_builer_inst(
			       .clock_and_control(),
			       .ttc_commands(),
			       .ctrl(),
			       .mon(),
			       .i_ptcalc(),
			       .i_pl2mtc(),
			       .o_mtc(),
			       .o_nsp()
			       );
   */
endmodule // end TopLevel module definition
