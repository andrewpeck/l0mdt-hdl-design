--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: rpc_z to tube windows 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library heg_roi_lib;
use heg_roi_lib.roi_types_pkg.all;

package RoI_LUT_BILA3 is

  constant BILA3_IN_MAX : integer := 540;

  -- type trLUT_limits_t is array (0 to 1) of integer;
  -- type trLUT_layer_t is array (0 to 5) of trLUT_limits_t; -- 1 layer has up to 212 z position
  -- type trLUT_station_t is array (0 to BILA3_IN_MAX) of trLUT_layer_t; -- 1 station has up to 6 layers
  -- type trLut_sector_t is array ( 0 to 3) of trLUT_station_t; -- 1 sector has 4 station

  constant trLUT_s3i_rom_mem : roi_mdt_lut := (
    0 to 240 => ((-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1)),  
    241 to 270 => ((-1,-1),(-1,-1),(-1,-1),(0,0),(0,0),(0,0)),  
    271 to 300 => ((0,0),(0,0),(0,0),(0,1),(0,1),(0,1)),  
    301 to 330 => ((0,1),(0,1),(0,1),(0,2),(0,2),(0,2)),  
    331 to 360 => ((0,2),(0,2),(0,2),(0,3),(0,3),(0,3)),  
    361 to 390 => ((0,3),(0,3),(0,3),(0,4),(0,4),(0,4)),  
    391 to 420 => ((0,4),(0,4),(0,4),(0,5),(0,5),(0,5)),  
    421 to 450 => ((0,5),(0,5),(0,5),(0,6),(0,6),(0,6)),  
    451 to 480 => ((0,6),(0,6),(0,6),(1,7),(1,7),(1,7)),  
    481 to 510 => ((1,7),(1,7),(1,7),(2,8),(2,8),(2,8)),  
    511 to 540 => ((2,8),(2,8),(2,8),(3,9),(3,9),(3,9)),
    541 to 1023 => ((0,0),(0,0),(0,0),(0,0),(0,0),(0,0))
  );

  --  constant trLUT_s3i_rom_mem : roi_mdt_lut := (
  --   0 to 240 => ((-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1)),  
  --   241 to 270 => ((-1,-1),(-1,-1),(-1,-1),(0,0),(0,0),(0,0)),  
  --   271 to 300 => ((0,0),(0,0),(0,0),(0,1),(0,1),(0,1)),  
  --   301 to 330 => ((0,1),(0,1),(0,1),(0,2),(0,2),(0,2)),  
  --   331 to 360 => ((0,2),(0,2),(0,2),(0,3),(0,3),(0,3)),  
  --   361 to 390 => ((0,3),(0,3),(0,3),(0,4),(0,4),(0,4)),  
  --   391 to 420 => ((0,4),(0,4),(0,4),(0,5),(0,5),(0,5)),  
  --   421 to 450 => ((0,5),(0,5),(0,5),(0,6),(0,6),(0,6)),  
  --   451 to 480 => ((0,6),(0,6),(0,6),(1,7),(1,7),(1,7)),  
  --   481 to 510 => ((1,7),(1,7),(1,7),(2,8),(2,8),(2,8)),  
  --   511 to 540 => ((2,8),(2,8),(2,8),(3,9),(3,9),(3,9)),
  --   541 to 1023 => ((0,0),(0,0),(0,0),(0,0),(0,0),(0,0))
  -- );

  -- constant trLUT_s3i_rom_mem : roi_mdt_lut := (
  --   0 to 240 => ((-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1)),  
  --   241 to 270 => ((-1,-1),(-1,-1),(-1,-1),(0,0),(0,0),(0,0)),  
  --   271 to 300 => ((0,0),(0,0),(0,0),(0,1),(0,1),(0,1)),  
  --   301 to 330 => ((0,1),(0,1),(0,1),(0,2),(0,2),(0,2)),  
  --   331 to 360 => ((0,2),(0,2),(0,2),(0,3),(0,3),(0,3)),  
  --   361 to 390 => ((0,3),(0,3),(0,3),(0,4),(0,4),(0,4)),  
  --   391 to 420 => ((0,4),(0,4),(0,4),(0,5),(0,5),(0,5)),  
  --   421 to 450 => ((0,5),(0,5),(0,5),(0,6),(0,6),(0,6)),  
  --   451 to 480 => ((0,6),(0,6),(0,6),(1,7),(1,7),(1,7)),  
  --   481 to 510 => ((1,7),(1,7),(1,7),(2,8),(2,8),(2,8)),  
  --   511 to 540 => ((2,8),(2,8),(2,8),(3,9),(3,9),(3,9)),  
  --   541 to 570 => ((3,9),(3,9),(3,9),(4,10),(4,10),(4,10)),  
  --   571 to 600 => ((4,10),(4,10),(4,10),(5,11),(5,11),(5,11)),  
  --   601 to 630 => ((4,10),(5,11),(5,11),(6,12),(6,12),(7,13)),  
  --   631 to 660 => ((5,11),(6,12),(6,12),(7,13),(7,13),(8,14)),  
  --   661 to 690 => ((6,12),(7,13),(7,13),(8,14),(9,15),(9,15)),  
  --   691 to 720 => ((7,13),(7,13),(8,14),(9,15),(10,16),(10,16)),  
  --   721 to 750 => ((8,14),(8,14),(9,15),(10,16),(11,17),(11,17)),  
  --   751 to 780 => ((9,15),(9,15),(10,16),(11,17),(12,18),(12,18)),  
  --   781 to 810 => ((10,16),(10,16),(11,17),(13,19),(13,19),(13,19)),  
  --   811 to 840 => ((11,17),(11,17),(11,17),(14,20),(14,20),(14,20)),  
  --   841 to 870 => ((12,18),(12,18),(12,18),(15,21),(15,21),(15,21)),  
  --   871 to 900 => ((13,19),(13,19),(13,19),(16,22),(16,22),(16,22)),  
  --   901 to 930 => ((14,20),(14,20),(14,20),(17,23),(17,23),(17,23)),  
  --   931 to 960 => ((15,21),(15,21),(15,21),(18,24),(18,24),(18,24)),  
  --   961 to 990 => ((16,22),(16,22),(16,22),(19,25),(19,25),(19,25)),  
  --   991 to 1020 => ((17,23),(17,23),(17,23),(20,26),(20,26),(20,26)),  
  --   1021 to 1050 => ((18,24),(18,24),(18,24),(21,27),(21,27),(21,27)),  
  --   1051 to 1080 => ((19,25),(19,25),(19,25),(22,28),(22,28),(22,28)),  
  --   1081 to 1110 => ((20,26),(20,26),(20,26),(23,29),(23,29),(23,29)),  
  --   1111 to 1140 => ((21,27),(21,27),(21,27),(24,30),(24,30),(24,30)),  
  --   1141 to 1170 => ((22,28),(22,28),(22,28),(25,30),(25,31),(25,31)),  
  --   1171 to 1200 => ((23,29),(23,29),(23,29),(26,31),(26,32),(27,32)),  
  --   1201 to 1230 => ((23,29),(24,30),(24,30),(27,32),(27,33),(28,33)),  
  --   1231 to 1260 => ((24,30),(25,30),(25,30),(28,33),(28,34),(29,34)),  
  --   1261 to 1290 => ((25,31),(26,31),(26,31),(29,34),(29,35),(30,35)),  
  --   1291 to 1320 => ((26,32),(27,32),(27,32),(30,36),(30,36),(30,36)),  
  --   1321 to 1350 => ((27,33),(28,33),(28,33),(31,37),(31,37),(31,37)),  
  --   1351 to 1380 => ((28,34),(28,34),(29,34),(32,38),(32,38),(32,38)),  
  --   1381 to 1410 => ((29,34),(29,35),(30,35),(33,39),(33,39),(33,39)),  
  --   1411 to 1440 => ((30,35),(30,36),(30,36),(34,40),(34,40),(34,40)),  
  --   1441 to 1470 => ((30,36),(31,37),(31,37),(35,41),(35,41),(35,41)),  
  --   1471 to 1500 => ((31,37),(32,38),(32,38),(36,42),(36,42),(36,42)),  
  --   1501 to 1530 => ((32,38),(33,39),(33,39),(37,43),(37,43),(37,43)),  
  --   1531 to 1560 => ((33,39),(34,40),(34,40),(38,44),(38,44),(38,44)),  
  --   1561 to 1590 => ((34,40),(34,40),(35,41),(39,45),(39,45),(40,46)),  
  --   1591 to 1620 => ((35,41),(35,41),(36,42),(40,46),(40,46),(41,47)),  
  --   1621 to 1650 => ((36,42),(36,42),(37,43),(41,47),(41,47),(42,48)),  
  --   1651 to 1680 => ((37,43),(37,43),(38,44),(42,48),(42,48),(43,49)),  
  --   1681 to 1710 => ((38,44),(38,44),(39,45),(43,49),(43,49),(44,50)),  
  --   1711 to 1740 => ((39,45),(39,45),(40,46),(44,50),(44,50),(45,51)),  
  --   1741 to 1770 => ((40,46),(40,46),(41,47),(45,51),(45,51),(46,52)),  
  --   1771 to 1800 => ((41,47),(41,47),(42,48),(46,52),(47,53),(47,53)),  
  --   1801 to 1830 => ((42,48),(42,48),(43,49),(47,53),(48,54),(48,54)),  
  --   1831 to 1860 => ((43,49),(43,49),(43,49),(48,54),(49,55),(49,55)),  
  --   1861 to 1890 => ((44,50),(44,50),(44,50),(49,55),(50,56),(50,56)),  
  --   1891 to 1920 => ((45,51),(45,51),(45,51),(50,56),(51,57),(51,57)),  
  --   1921 to 1950 => ((46,52),(46,52),(46,52),(51,57),(52,58),(52,58)),  
  --   1951 to 1980 => ((47,53),(47,53),(47,53),(52,58),(53,59),(53,59)),  
  --   1981 to 2010 => ((47,53),(48,54),(48,54),(53,59),(54,60),(54,60)),  
  --   2011 to 2040 => ((48,54),(49,55),(49,55),(54,60),(55,61),(55,61)),  
  --   2041 to 2070 => ((49,55),(50,56),(50,56),(56,62),(56,62),(56,62)),  
  --   2071 to 2100 => ((50,56),(51,57),(51,57),(57,63),(57,63),(57,63)),  
  --   2101 to 2130 => ((51,57),(52,58),(52,58),(58,64),(58,64),(58,64)),  
  --   2131 to 2160 => ((52,58),(53,59),(53,59),(59,65),(59,65),(60,66)),  
  --   2161 to 2190 => ((53,59),(54,60),(54,60),(60,66),(60,66),(61,66)),  
  --   2191 to 2220 => ((54,60),(55,61),(55,61),(61,66),(61,66),(62,67)),  
  --   2221 to 2250 => ((55,61),(56,62),(56,62),(62,67),(62,68),(63,68)),  
  --   2251 to 2280 => ((56,62),(56,62),(57,63),(63,68),(63,69),(64,69)),  
  --   2281 to 2310 => ((57,63),(57,63),(58,64),(64,69),(64,70),(65,70)),  
  --   2311 to 2340 => ((58,64),(58,64),(59,65),(65,70),(65,71),(66,71)),  
  --   2341 to 2370 => ((59,65),(59,65),(60,66),(66,71),(66,72),(66,72)),  
  --   2371 to 2400 => ((60,66),(60,66),(61,66),(66,72),(67,73),(67,73)),  
  --   2401 to 2430 => ((61,66),(61,67),(62,67),(67,73),(68,74),(68,74)),  
  --   2431 to 2460 => ((62,67),(62,68),(63,68),(68,74),(69,75),(69,75)),  
  --   2461 to 2490 => ((63,68),(63,68),(64,69),(69,75),(70,76),(70,76)),  
  --   2491 to 2520 => ((64,69),(64,69),(65,70),(70,76),(71,77),(71,77)),  
  --   2521 to 2550 => ((65,70),(65,70),(66,71),(71,77),(72,78),(73,79)),  
  --   2551 to 2580 => ((65,71),(66,71),(66,72),(72,78),(73,79),(74,80)),  
  --   2581 to 2610 => ((66,72),(66,72),(67,73),(74,80),(74,80),(75,81)),  
  --   2611 to 2640 => ((67,73),(67,73),(68,74),(75,81),(75,81),(76,82)),  
  --   2641 to 2670 => ((68,74),(68,74),(69,75),(76,82),(76,82),(77,83)),  
  --   2671 to 2700 => ((69,75),(69,75),(70,76),(77,83),(77,83),(78,84)),  
  --   2701 to 2730 => ((70,76),(70,76),(71,77),(78,84),(78,84),(79,85)),  
  --   2731 to 2760 => ((70,76),(71,77),(72,78),(79,85),(79,85),(80,86)),  
  --   2761 to 2790 => ((71,77),(72,78),(73,79),(80,86),(80,86),(81,87)),  
  --   2791 to 2820 => ((72,78),(73,79),(74,80),(81,87),(81,87),(82,88)),  
  --   2821 to 2850 => ((73,79),(74,80),(75,81),(82,88),(82,88),(83,89)),  
  --   2851 to 2880 => ((74,80),(75,81),(75,81),(83,89),(83,89),(84,90)),  
  --   2881 to 2910 => ((75,81),(76,82),(76,82),(84,90),(85,91),(85,91)),  
  --   2911 to 2940 => ((76,82),(77,83),(77,83),(85,91),(86,92),(86,92)),  
  --   2941 to 2970 => ((77,83),(78,84),(78,84),(86,92),(87,93),(87,93)),  
  --   2971 to 3000 => ((78,84),(79,85),(79,85),(87,93),(88,94),(88,94)),  
  --   3001 to 3030 => ((79,85),(80,86),(80,86),(88,94),(89,95),(89,95)),  
  --   3031 to 3060 => ((80,86),(81,87),(81,87),(89,95),(90,96),(90,96)),  
  --   3061 to 3090 => ((81,87),(82,88),(82,88),(90,96),(91,97),(91,97)),  
  --   3091 to 3120 => ((82,88),(83,89),(83,89),(91,97),(92,98),(93,99)),  
  --   3121 to 3150 => ((83,89),(83,89),(84,90),(92,98),(93,99),(94,100)),  
  --   3151 to 3180 => ((84,90),(84,90),(85,91),(93,99),(94,100),(95,101)),  
  --   3181 to 3210 => ((85,91),(85,91),(86,92),(94,100),(95,101),(96,102)),  
  --   3211 to 3240 => ((86,92),(86,92),(87,93),(95,101),(96,102),(97,96)),  
  --   3241 to 3270 => ((87,93),(87,93),(88,94),(96,96),(97,96),(98,97)),  
  --   3271 to 3300 => ((88,94),(88,94),(89,95),(97,97),(98,97),(99,98)),  
  --   3301 to 3330 => ((89,95),(89,95),(90,96),(98,98),(99,98),(100,99)),  
  --   3331 to 3360 => ((89,95),(90,96),(91,97),(100,99),(100,100),(101,100)),  
  --   3361 to 3390 => ((90,96),(91,97),(92,98),(101,100),(101,101),(102,101)),  
  --   3391 to 3420 => ((91,97),(92,98),(93,99),(102,101),(96,102),(96,102)),  
  --   3421 to 3450 => ((92,98),(93,99),(94,100),(96,102),(97,103),(97,103)),  
  --   3451 to 3480 => ((93,99),(94,100),(95,101),(97,103),(98,104),(98,104)),  
  --   3481 to 3510 => ((94,100),(95,101),(96,102),(98,104),(99,105),(99,105)),  
  --   3511 to 3540 => ((95,101),(96,102),(97,96),(99,105),(100,106),(101,107)),  
  --   3541 to 3570 => ((96,102),(97,96),(98,97),(100,106),(101,107),(102,108)),  
  --   3571 to 3600 => ((97,96),(98,97),(99,98),(101,107),(102,108),(103,109)),  
  --   3601 to 3630 => ((98,97),(99,98),(100,99),(102,108),(103,109),(104,110)),  
  --   3631 to 3660 => ((99,98),(100,99),(100,100),(103,109),(104,110),(105,111)),  
  --   3661 to 3690 => ((100,99),(101,100),(101,101),(104,110),(105,111),(106,112)),  
  --   3691 to 3720 => ((101,100),(102,101),(96,102),(105,111),(106,112),(107,113)),  
  --   3721 to 3750 => ((102,101),(96,102),(97,103),(106,112),(107,113),(108,114)),  
  --   3751 to 3780 => ((96,102),(97,103),(98,104),(107,113),(108,114),(109,115)),  
  --   3781 to 3810 => ((97,103),(98,104),(99,105),(108,114),(109,115),(110,116)),  
  --   3811 to 3840 => ((98,104),(99,105),(100,106),(109,115),(110,116),(111,117)),  
  --   3841 to 3870 => ((99,105),(100,106),(101,107),(110,116),(111,117),(112,118)),  
  --   3871 to 3900 => ((100,106),(101,107),(101,107),(112,118),(112,118),(113,119)),  
  --   3901 to 3930 => ((101,107),(102,108),(102,108),(113,119),(113,119),(114,120)),  
  --   3931 to 3960 => ((102,108),(103,109),(103,109),(114,120),(114,120),(115,121)),  
  --   3961 to 3990 => ((103,109),(104,110),(104,110),(115,121),(115,121),(116,122)),  
  --   3991 to 4020 => ((104,110),(105,111),(105,111),(116,122),(117,123),(117,123)),  
  --   4021 to 4050 => ((105,111),(105,111),(106,112),(117,123),(118,124),(118,124)),  
  --   4051 to 4080 => ((106,112),(106,112),(107,113),(118,124),(119,125),(119,125)),  
  --   4081 to 4110 => ((107,113),(107,113),(108,114),(119,125),(120,126),(121,127)),  
  --   4111 to 4140 => ((107,113),(108,114),(109,115),(120,126),(121,127),(122,128)),  
  --   4141 to 4170 => ((108,114),(109,115),(110,116),(121,127),(122,128),(123,129)),  
  --   4171 to 4200 => ((109,115),(110,116),(111,117),(122,128),(123,129),(124,130)),  
  --   4201 to 4230 => ((110,116),(111,117),(112,118),(123,129),(124,130),(125,131)),  
  --   4231 to 4260 => ((111,117),(112,118),(113,119),(124,130),(125,131),(126,132)),  
  --   4261 to 4290 => ((112,118),(113,119),(114,120),(125,131),(126,132),(127,132)),  
  --   4291 to 4320 => ((113,119),(114,120),(115,121),(126,132),(127,132),(128,133)),  
  --   4321 to 4350 => ((114,120),(115,121),(116,122),(127,132),(128,133),(129,134)),  
  --   4351 to 4380 => ((115,121),(116,122),(117,123),(128,133),(129,134),(130,135)),  
  --   4381 to 4410 => ((116,122),(117,123),(118,124),(129,135),(130,135),(131,136)),  
  --   4411 to 4440 => ((117,123),(118,124),(119,125),(130,136),(131,136),(132,137)),  
  --   4441 to 4470 => ((118,124),(119,125),(120,126),(131,137),(132,138),(132,138)),  
  --   4471 to 4500 => ((119,125),(120,126),(121,127),(132,138),(133,139),(134,140)),  
  --   4501 to 4530 => ((120,126),(121,127),(122,128),(133,139),(134,140),(135,141)),  
  --   4531 to 4560 => ((121,127),(122,128),(123,129),(134,140),(135,141),(136,142)),  
  --   4561 to 4590 => ((122,128),(123,129),(124,130),(135,141),(136,142),(137,143)),  
  --   4591 to 4620 => ((123,129),(124,130),(125,131),(136,142),(137,143),(138,144)),  
  --   4621 to 4650 => ((124,130),(125,131),(126,132),(137,143),(138,144),(139,145)),  
  --   4651 to 4680 => ((125,131),(126,132),(127,132),(138,144),(139,145),(140,146)),  
  --   4681 to 4710 => ((125,131),(126,132),(127,133),(139,145),(140,146),(141,147)),  
  --   4711 to 4740 => ((126,132),(127,133),(128,134),(140,146),(141,147),(142,148)),  
  --   4741 to 4770 => ((127,133),(128,134),(129,135),(141,147),(142,148),(143,149)),  
  --   4771 to 4800 => ((128,134),(129,135),(130,136),(142,148),(143,149),(144,150)),  
  --   4801 to 4830 => ((129,135),(130,136),(131,137),(143,149),(144,150),(145,151)),  
  --   4831 to 4860 => ((130,136),(131,137),(132,138),(144,150),(145,151),(146,152)),  
  --   4861 to 4890 => ((131,136),(132,138),(133,139),(145,151),(146,152),(147,153)),  
  --   4891 to 4920 => ((132,137),(132,138),(133,139),(146,152),(147,153),(148,154)),  
  --   4921 to 4950 => ((132,138),(133,139),(134,140),(147,153),(148,154),(149,155)),  
  --   4951 to 4980 => ((133,139),(134,140),(135,141),(148,154),(149,155),(150,156)),  
  --   4981 to 5010 => ((134,140),(135,141),(136,142),(149,155),(150,156),(151,157)),  
  --   5011 to 5040 => ((135,141),(136,142),(137,143),(150,156),(151,157),(152,158)),  
  --   5041 to 5070 => ((136,142),(137,143),(138,144),(151,157),(152,158),(154,160)),  
  --   5071 to 5100 => ((137,143),(138,144),(139,145),(152,158),(153,159),(155,161)),  
  --   5101 to 5130 => ((138,144),(139,145),(140,146),(153,159),(155,161),(156,162)),  
  --   5131 to 5160 => ((139,145),(140,146),(141,147),(155,161),(156,162),(157,162)),  
  --   5161 to 5190 => ((140,146),(141,147),(142,148),(156,162),(157,162),(158,163)),  
  --   5191 to 5220 => ((141,147),(142,148),(143,149),(157,162),(158,163),(159,164)),  
  --   5221 to 5250 => ((142,148),(143,149),(144,150),(158,163),(159,164),(160,165)),  
  --   5251 to 5280 => ((143,149),(144,150),(145,151),(159,164),(160,165),(161,166)),  
  --   5281 to 5310 => ((144,150),(145,151),(146,152),(160,165),(161,166),(162,167)),  
  --   5311 to 5340 => ((145,151),(146,152),(147,153),(161,166),(162,167),(162,168)),  
  --   5341 to 5370 => ((146,152),(147,153),(148,154),(162,167),(162,168),(163,169)),  
  --   5371 to 5400 => ((147,153),(148,154),(149,155),(162,168),(163,169),(164,170)),  
  --   5401 to 5430 => ((148,154),(149,155),(150,156),(163,169),(164,170),(165,171)),  
  --   5431 to 5460 => ((149,155),(150,156),(151,157),(164,170),(165,171),(166,172)),  
  --   5461 to 5490 => ((149,155),(151,157),(152,158),(165,171),(166,172),(168,174)),  
  --   5491 to 5520 => ((150,156),(152,158),(153,159),(166,172),(167,173),(169,175)),  
  --   5521 to 5550 => ((151,157),(153,159),(154,160),(167,173),(168,174),(170,176)),  
  --   5551 to 5580 => ((152,158),(153,159),(155,161),(168,174),(170,176),(171,177)),  
  --   5581 to 5610 => ((153,159),(154,160),(156,162),(169,175),(171,177),(172,178)),  
  --   5611 to 5640 => ((154,160),(155,161),(157,162),(170,176),(172,178),(173,179)),  
  --   5641 to 5670 => ((155,161),(156,162),(158,163),(171,177),(173,179),(174,180)),  
  --   5671 to 5700 => ((156,162),(157,163),(159,164),(173,179),(174,180),(175,181)),  
  --   5701 to 5730 => ((157,162),(158,164),(159,165),(174,180),(175,181),(176,182)),  
  --   5731 to 5760 => ((158,163),(159,165),(160,166),(175,181),(176,182),(177,183)),  
  --   5761 to 5790 => ((159,164),(160,165),(161,167),(176,182),(177,183),(178,184)),  
  --   5791 to 5820 => ((160,165),(161,166),(162,168),(177,183),(178,184),(179,185)),  
  --   5821 to 5850 => ((161,166),(162,167),(163,169),(178,184),(179,185),(180,186)),  
  --   5851 to 5880 => ((162,167),(162,168),(164,170),(179,185),(180,186),(181,187)),  
  --   5881 to 5910 => ((162,168),(163,169),(165,171),(180,186),(181,187),(182,188)),  
  --   5911 to 5940 => ((163,169),(164,170),(166,172),(181,187),(182,188),(183,189)),  
  --   5941 to 5970 => ((164,170),(165,171),(166,172),(182,188),(183,189),(184,190)),  
  --   5971 to 6000 => ((165,171),(166,172),(167,173),(183,189),(184,190),(185,191)),  
  --   6001 to 6030 => ((166,172),(167,173),(168,174),(184,190),(185,191),(186,192)),  
  --   6031 to 6060 => ((167,173),(168,174),(169,175),(185,191),(186,192),(188,194)),  
  --   6061 to 6090 => ((168,174),(169,175),(170,176),(186,192),(187,193),(189,195)),  
  --   6091 to 6120 => ((169,175),(170,176),(171,177),(187,193),(188,194),(190,196)),  
  --   6121 to 6150 => ((170,176),(171,177),(172,178),(188,194),(189,195),(191,197)),  
  --   6151 to 6180 => ((171,177),(172,178),(173,179),(189,195),(190,196),(192,198)),  
  --   6181 to 6210 => ((172,178),(173,179),(174,180),(190,196),(192,198),(193,199)),  
  --   6211 to 6240 => ((173,179),(174,180),(175,181),(191,197),(193,199),(194,200)),  
  --   6241 to 6270 => ((173,179),(175,181),(176,182),(192,198),(194,200),(195,201)),  
  --   6271 to 6300 => ((174,180),(176,182),(177,183),(193,199),(195,201),(196,202)),  
  --   6301 to 6330 => ((175,181),(177,183),(178,184),(194,200),(196,202),(197,203)),  
  --   6331 to 6360 => ((176,182),(178,184),(179,185),(195,201),(197,203),(198,204)),  
  --   6361 to 6390 => ((177,183),(179,185),(180,186),(196,202),(198,204),(199,205)),  
  --   6391 to 6420 => ((178,184),(180,186),(181,187),(197,203),(199,205),(200,206)),  
  --   6421 to 6450 => ((179,185),(181,187),(182,188),(199,205),(200,206),(201,207)),  
  --   6451 to 6480 => ((180,186),(181,187),(183,189),(200,206),(201,207),(202,208)),  
  --   6481 to 6510 => ((181,187),(182,188),(184,190),(201,207),(202,208),(203,209)),  
  --   6511 to 6550 => ((182,188),(183,189),(185,191),(202,208),(203,209),(204,210)),
  --   6551 to 13000 => ((0,0),(0,0),(0,0),(0,0),(0,0),(0,0))
  -- );

 end package RoI_LUT_BILA3;
