

 get_rom_addr get_rom_addr_inst(
	       .ap_clk(clk),
	       .ap_rst(ap_rst_gra), //|hba_reset_fo[0]),
	       .ap_start(gra_ap_start),
	       .ap_done(gra_ap_done),
	       .ap_idle(gra_ap_idle),
	       .ap_ready(gra_ap_ready),
	       .in_val_V_ap_vld(gra_theta_vld),
	       .in_val_V(gra_theta),
				.total_bins_V(gra_total_bins),
	       .sin_rom_addr_0_V(sin_rom_addr_start[0]),
	       .sin_rom_addr_0_V_ap_vld(),
	       .sin_rom_addr_1_V(sin_rom_addr_start[1]),
	       .sin_rom_addr_1_V_ap_vld(),
	       .sin_rom_addr_2_V(sin_rom_addr_start[2]),
	       .sin_rom_addr_2_V_ap_vld(),
	       .sin_rom_addr_3_V(sin_rom_addr_start[3]),
	       .sin_rom_addr_3_V_ap_vld(),
	       .sin_rom_addr_4_V(sin_rom_addr_start[4]),
	       .sin_rom_addr_4_V_ap_vld(),
	       .sin_rom_addr_5_V(sin_rom_addr_start[5]),
	       .sin_rom_addr_5_V_ap_vld(),
	       .sin_rom_addr_6_V(sin_rom_addr_start[6]),
	       .sin_rom_addr_6_V_ap_vld(),
	       .sin_rom_addr_7_V(sin_rom_addr_start[7]),
	       .sin_rom_addr_7_V_ap_vld(),
	       .sin_rom_addr_8_V(sin_rom_addr_start[8]),
	       .sin_rom_addr_8_V_ap_vld(),
	       .sin_rom_addr_9_V(sin_rom_addr_start[9]),
	       .sin_rom_addr_9_V_ap_vld(),
	       .sin_rom_addr_10_V(sin_rom_addr_start[10]),
	       .sin_rom_addr_10_V_ap_vld(),
	       .sin_rom_addr_11_V(sin_rom_addr_start[11]),
	       .sin_rom_addr_11_V_ap_vld(),
	       .sin_rom_addr_12_V(sin_rom_addr_start[12]),
	       .sin_rom_addr_12_V_ap_vld(),
	       .sin_rom_addr_13_V(sin_rom_addr_start[13]),
	       .sin_rom_addr_13_V_ap_vld(),
	       .sin_rom_addr_14_V(sin_rom_addr_start[14]),
	       .sin_rom_addr_14_V_ap_vld(),
	       .sin_rom_addr_15_V(sin_rom_addr_start[15]),
	       .sin_rom_addr_15_V_ap_vld(),
	       .sin_rom_sel_0_V(sin_rom_sel[0]),
	       .sin_rom_sel_0_V_ap_vld(),
	       .sin_rom_sel_1_V(sin_rom_sel[1]),
	       .sin_rom_sel_1_V_ap_vld(),
	       .sin_rom_sel_2_V(sin_rom_sel[2]),
	       .sin_rom_sel_2_V_ap_vld(),
	       .sin_rom_sel_3_V(sin_rom_sel[3]),
	       .sin_rom_sel_3_V_ap_vld(),
	       .sin_rom_sel_4_V(sin_rom_sel[4]),
	       .sin_rom_sel_4_V_ap_vld(),
	       .sin_rom_sel_5_V(sin_rom_sel[5]),
	       .sin_rom_sel_5_V_ap_vld(),
	       .sin_rom_sel_6_V(sin_rom_sel[6]),
	       .sin_rom_sel_6_V_ap_vld(),
	       .sin_rom_sel_7_V(sin_rom_sel[7]),
	       .sin_rom_sel_7_V_ap_vld(),
	       .sin_rom_sel_8_V(sin_rom_sel[8]),
	       .sin_rom_sel_8_V_ap_vld(),
	       .sin_rom_sel_9_V(sin_rom_sel[9]),
	       .sin_rom_sel_9_V_ap_vld(),
	       .sin_rom_sel_10_V(sin_rom_sel[10]),
	       .sin_rom_sel_10_V_ap_vld(),
	       .sin_rom_sel_11_V(sin_rom_sel[11]),
	       .sin_rom_sel_11_V_ap_vld(),
	       .sin_rom_sel_12_V(sin_rom_sel[12]),
	       .sin_rom_sel_12_V_ap_vld(),
	       .sin_rom_sel_13_V(sin_rom_sel[13]),
	       .sin_rom_sel_13_V_ap_vld(),
	       .sin_rom_sel_14_V(sin_rom_sel[14]),
	       .sin_rom_sel_14_V_ap_vld(),
	       .sin_rom_sel_15_V(sin_rom_sel[15]),
	       .sin_rom_sel_15_V_ap_vld(),
	       .cos_rom_addr_0_V(cos_rom_addr_start[0]),
	       .cos_rom_addr_0_V_ap_vld(),
	       .cos_rom_addr_1_V(cos_rom_addr_start[1]),
	       .cos_rom_addr_1_V_ap_vld(),
	       .cos_rom_addr_2_V(cos_rom_addr_start[2]),
	       .cos_rom_addr_2_V_ap_vld(),
	       .cos_rom_addr_3_V(cos_rom_addr_start[3]),
	       .cos_rom_addr_3_V_ap_vld(),
	       .cos_rom_addr_4_V(cos_rom_addr_start[4]),
	       .cos_rom_addr_4_V_ap_vld(),
	       .cos_rom_addr_5_V(cos_rom_addr_start[5]),
	       .cos_rom_addr_5_V_ap_vld(),
	       .cos_rom_addr_6_V(cos_rom_addr_start[6]),
	       .cos_rom_addr_6_V_ap_vld(),
	       .cos_rom_addr_7_V(cos_rom_addr_start[7]),
	       .cos_rom_addr_7_V_ap_vld(),
	       .cos_rom_addr_8_V(cos_rom_addr_start[8]),
	       .cos_rom_addr_8_V_ap_vld(),
	       .cos_rom_addr_9_V(cos_rom_addr_start[9]),
	       .cos_rom_addr_9_V_ap_vld(),
	       .cos_rom_addr_10_V(cos_rom_addr_start[10]),
	       .cos_rom_addr_10_V_ap_vld(),
	       .cos_rom_addr_11_V(cos_rom_addr_start[11]),
	       .cos_rom_addr_11_V_ap_vld(),
	       .cos_rom_addr_12_V(cos_rom_addr_start[12]),
	       .cos_rom_addr_12_V_ap_vld(),
	       .cos_rom_addr_13_V(cos_rom_addr_start[13]),
	       .cos_rom_addr_13_V_ap_vld(),
	       .cos_rom_addr_14_V(cos_rom_addr_start[14]),
	       .cos_rom_addr_14_V_ap_vld(),
	       .cos_rom_addr_15_V(cos_rom_addr_start[15]),
	       .cos_rom_addr_15_V_ap_vld(),
	       .cos_rom_sel_0_V(cos_rom_sel[0]),
	       .cos_rom_sel_0_V_ap_vld(),
	       .cos_rom_sel_1_V(cos_rom_sel[1]),
	       .cos_rom_sel_1_V_ap_vld(),
	       .cos_rom_sel_2_V(cos_rom_sel[2]),
	       .cos_rom_sel_2_V_ap_vld(),
	       .cos_rom_sel_3_V(cos_rom_sel[3]),
	       .cos_rom_sel_3_V_ap_vld(),
	       .cos_rom_sel_4_V(cos_rom_sel[4]),
	       .cos_rom_sel_4_V_ap_vld(),
	       .cos_rom_sel_5_V(cos_rom_sel[5]),
	       .cos_rom_sel_5_V_ap_vld(),
	       .cos_rom_sel_6_V(cos_rom_sel[6]),
	       .cos_rom_sel_6_V_ap_vld(),
	       .cos_rom_sel_7_V(cos_rom_sel[7]),
	       .cos_rom_sel_7_V_ap_vld(),
	       .cos_rom_sel_8_V(cos_rom_sel[8]),
	       .cos_rom_sel_8_V_ap_vld(),
	       .cos_rom_sel_9_V(cos_rom_sel[9]),
	       .cos_rom_sel_9_V_ap_vld(),
	       .cos_rom_sel_10_V(cos_rom_sel[10]),
	       .cos_rom_sel_10_V_ap_vld(),
	       .cos_rom_sel_11_V(cos_rom_sel[11]),
	       .cos_rom_sel_11_V_ap_vld(),
	       .cos_rom_sel_12_V(cos_rom_sel[12]),
	       .cos_rom_sel_12_V_ap_vld(),
	       .cos_rom_sel_13_V(cos_rom_sel[13]),
	       .cos_rom_sel_13_V_ap_vld(),
	       .cos_rom_sel_14_V(cos_rom_sel[14]),
	       .cos_rom_sel_14_V_ap_vld(),
	       .cos_rom_sel_15_V(cos_rom_sel[15]),
	       .cos_rom_sel_15_V_ap_vld()
	       );


get_trig_vals get_trig_vals_inst(
				 .ap_clk(clk),
				 .ap_rst((ap_rst_gra)), // | hba_reset)),
				 .ap_start(get_next_rom_addr),//theta_offset_factor_sn_vld_128),//sin_addr_offset_V_TVALID),
				 .ap_done(gtv_ap_done),
				 .ap_idle(gtv_ap_idle),
				 .ap_ready(gtv_ap_ready),
				 .sin_addr_base_0_V(sin_rom_addr[0]),
				 .sin_addr_base_1_V(sin_rom_addr[1]),
				 .sin_addr_base_2_V(sin_rom_addr[2]),
				 .sin_addr_base_3_V(sin_rom_addr[3]),
				 .sin_addr_base_4_V(sin_rom_addr[4]),
				 .sin_addr_base_5_V(sin_rom_addr[5]),
				 .sin_addr_base_6_V(sin_rom_addr[6]),
				 .sin_addr_base_7_V(sin_rom_addr[7]),
				 .sin_addr_base_8_V(sin_rom_addr[8]),
				 .sin_addr_base_9_V(sin_rom_addr[9]),
				 .sin_addr_base_10_V(sin_rom_addr[10]),
				 .sin_addr_base_11_V(sin_rom_addr[11]),
				 .sin_addr_base_12_V(sin_rom_addr[12]),
				 .sin_addr_base_13_V(sin_rom_addr[13]),
				 .sin_addr_base_14_V(sin_rom_addr[14]),
				 .sin_addr_base_15_V(sin_rom_addr[15]),
				 .hw_sin_val_8_0_V(hw_sin_val_16[0][23:16]),
				 .hw_sin_val_8_0_V_ap_vld(hw_sin_val_vld),
				 .hw_sin_val_8_1_V(hw_sin_val_16[1][23:16]),
				 .hw_sin_val_8_1_V_ap_vld(),
				 .hw_sin_val_8_2_V(hw_sin_val_16[2][23:16]),
				 .hw_sin_val_8_2_V_ap_vld(),
				 .hw_sin_val_8_3_V(hw_sin_val_16[3][23:16]),
				 .hw_sin_val_8_3_V_ap_vld(),
				 .hw_sin_val_8_4_V(hw_sin_val_16[4][23:16]),
				 .hw_sin_val_8_4_V_ap_vld(),
				 .hw_sin_val_8_5_V(hw_sin_val_16[5][23:16]),
				 .hw_sin_val_8_5_V_ap_vld(),
				 .hw_sin_val_8_6_V(hw_sin_val_16[6][23:16]),
				 .hw_sin_val_8_6_V_ap_vld(),
				 .hw_sin_val_8_7_V(hw_sin_val_16[7][23:16]),
				 .hw_sin_val_8_7_V_ap_vld(),
				 .hw_sin_val_8_8_V(hw_sin_val_16[8][23:16]),
				 .hw_sin_val_8_8_V_ap_vld(),
				 .hw_sin_val_8_9_V(hw_sin_val_16[9][23:16]),
				 .hw_sin_val_8_9_V_ap_vld(),
				 .hw_sin_val_8_10_V(hw_sin_val_16[10][23:16]),
				 .hw_sin_val_8_10_V_ap_vld(),
				 .hw_sin_val_8_11_V(hw_sin_val_16[11][23:16]),
				 .hw_sin_val_8_11_V_ap_vld(),
				 .hw_sin_val_8_12_V(hw_sin_val_16[12][23:16]),
				 .hw_sin_val_8_12_V_ap_vld(),
				 .hw_sin_val_8_13_V(hw_sin_val_16[13][23:16]),
				 .hw_sin_val_8_13_V_ap_vld(),
				 .hw_sin_val_8_14_V(hw_sin_val_16[14][23:16]),
				 .hw_sin_val_8_14_V_ap_vld(),
				 .hw_sin_val_8_15_V(hw_sin_val_16[15][23:16]),
				 .hw_sin_val_8_15_V_ap_vld(),
				 .hw_sin_val_16_0_V(hw_sin_val_16[0][15:0]),
				 .hw_sin_val_16_0_V_ap_vld(),
				 .hw_sin_val_16_1_V(hw_sin_val_16[1][15:0]),
				 .hw_sin_val_16_1_V_ap_vld(),
				 .hw_sin_val_16_2_V(hw_sin_val_16[2][15:0]),
				 .hw_sin_val_16_2_V_ap_vld(),
				 .hw_sin_val_16_3_V(hw_sin_val_16[3][15:0]),
				 .hw_sin_val_16_3_V_ap_vld(),
				 .hw_sin_val_16_4_V(hw_sin_val_16[4][15:0]),
				 .hw_sin_val_16_4_V_ap_vld(),
				 .hw_sin_val_16_5_V(hw_sin_val_16[5][15:0]),
				 .hw_sin_val_16_5_V_ap_vld(),
				 .hw_sin_val_16_6_V(hw_sin_val_16[6][15:0]),
				 .hw_sin_val_16_6_V_ap_vld(),
				 .hw_sin_val_16_7_V(hw_sin_val_16[7][15:0]),
				 .hw_sin_val_16_7_V_ap_vld(),
				 .hw_sin_val_16_8_V(hw_sin_val_16[8][15:0]),
				 .hw_sin_val_16_8_V_ap_vld(),
				 .hw_sin_val_16_9_V(hw_sin_val_16[9][15:0]),
				 .hw_sin_val_16_9_V_ap_vld(),
				 .hw_sin_val_16_10_V(hw_sin_val_16[10][15:0]),
				 .hw_sin_val_16_10_V_ap_vld(),
				 .hw_sin_val_16_11_V(hw_sin_val_16[11][15:0]),
				 .hw_sin_val_16_11_V_ap_vld(),
				 .hw_sin_val_16_12_V(hw_sin_val_16[12][15:0]),
				 .hw_sin_val_16_12_V_ap_vld(),
				 .hw_sin_val_16_13_V(hw_sin_val_16[13][15:0]),
				 .hw_sin_val_16_13_V_ap_vld(),
				 .hw_sin_val_16_14_V(hw_sin_val_16[14][15:0]),
				 .hw_sin_val_16_14_V_ap_vld(),
				 .hw_sin_val_16_15_V(hw_sin_val_16[15][15:0]),
				 .hw_sin_val_16_15_V_ap_vld(),
				 .sin_rom_sel_0_V(sin_rom_sel_reg[0]),
				 .sin_rom_sel_1_V(sin_rom_sel_reg[1]),
				 .sin_rom_sel_2_V(sin_rom_sel_reg[2]),
				 .sin_rom_sel_3_V(sin_rom_sel_reg[3]),
				 .sin_rom_sel_4_V(sin_rom_sel_reg[4]),
				 .sin_rom_sel_5_V(sin_rom_sel_reg[5]),
				 .sin_rom_sel_6_V(sin_rom_sel_reg[6]),
				 .sin_rom_sel_7_V(sin_rom_sel_reg[7]),
				 .sin_rom_sel_8_V(sin_rom_sel_reg[8]),
				 .sin_rom_sel_9_V(sin_rom_sel_reg[9]),
				 .sin_rom_sel_10_V(sin_rom_sel_reg[10]),
				 .sin_rom_sel_11_V(sin_rom_sel_reg[11]),
				 .sin_rom_sel_12_V(sin_rom_sel_reg[12]),
				 .sin_rom_sel_13_V(sin_rom_sel_reg[13]),
				 .sin_rom_sel_14_V(sin_rom_sel_reg[14]),
				 .sin_rom_sel_15_V(sin_rom_sel_reg[15]),
				 .cos_addr_base_0_V(cos_rom_addr[0]),
				 .cos_addr_base_1_V(cos_rom_addr[1]),
				 .cos_addr_base_2_V(cos_rom_addr[2]),
				 .cos_addr_base_3_V(cos_rom_addr[3]),
				 .cos_addr_base_4_V(cos_rom_addr[4]),
				 .cos_addr_base_5_V(cos_rom_addr[5]),
				 .cos_addr_base_6_V(cos_rom_addr[6]),
				 .cos_addr_base_7_V(cos_rom_addr[7]),
				 .cos_addr_base_8_V(cos_rom_addr[8]),
				 .cos_addr_base_9_V(cos_rom_addr[9]),
				 .cos_addr_base_10_V(cos_rom_addr[10]),
				 .cos_addr_base_11_V(cos_rom_addr[11]),
				 .cos_addr_base_12_V(cos_rom_addr[12]),
				 .cos_addr_base_13_V(cos_rom_addr[13]),
				 .cos_addr_base_14_V(cos_rom_addr[14]),
				 .cos_addr_base_15_V(cos_rom_addr[15]),
				 .hw_cos_val_8_0_V(hw_cos_val_16[0][23:16]),
				 .hw_cos_val_8_0_V_ap_vld(hw_cos_val_vld),
				 .hw_cos_val_8_1_V(hw_cos_val_16[1][23:16]),
				 .hw_cos_val_8_1_V_ap_vld(),
				 .hw_cos_val_8_2_V(hw_cos_val_16[2][23:16]),
				 .hw_cos_val_8_2_V_ap_vld(),
				 .hw_cos_val_8_3_V(hw_cos_val_16[3][23:16]),
				 .hw_cos_val_8_3_V_ap_vld(),
				 .hw_cos_val_8_4_V(hw_cos_val_16[4][23:16]),
				 .hw_cos_val_8_4_V_ap_vld(),
				 .hw_cos_val_8_5_V(hw_cos_val_16[5][23:16]),
				 .hw_cos_val_8_5_V_ap_vld(),
				 .hw_cos_val_8_6_V(hw_cos_val_16[6][23:16]),
				 .hw_cos_val_8_6_V_ap_vld(),
				 .hw_cos_val_8_7_V(hw_cos_val_16[7][23:16]),
				 .hw_cos_val_8_7_V_ap_vld(),
				 .hw_cos_val_8_8_V(hw_cos_val_16[8][23:16]),
				 .hw_cos_val_8_8_V_ap_vld(),
				 .hw_cos_val_8_9_V(hw_cos_val_16[9][23:16]),
				 .hw_cos_val_8_9_V_ap_vld(),
				 .hw_cos_val_8_10_V(hw_cos_val_16[10][23:16]),
				 .hw_cos_val_8_10_V_ap_vld(),
				 .hw_cos_val_8_11_V(hw_cos_val_16[11][23:16]),
				 .hw_cos_val_8_11_V_ap_vld(),
				 .hw_cos_val_8_12_V(hw_cos_val_16[12][23:16]),
				 .hw_cos_val_8_12_V_ap_vld(),
				 .hw_cos_val_8_13_V(hw_cos_val_16[13][23:16]),
				 .hw_cos_val_8_13_V_ap_vld(),
				 .hw_cos_val_8_14_V(hw_cos_val_16[14][23:16]),
				 .hw_cos_val_8_14_V_ap_vld(),
				 .hw_cos_val_8_15_V(hw_cos_val_16[15][23:16]),
				 .hw_cos_val_8_15_V_ap_vld(),
				 .hw_cos_val_16_0_V(hw_cos_val_16[0][15:0]),
				 .hw_cos_val_16_0_V_ap_vld(),
				 .hw_cos_val_16_1_V(hw_cos_val_16[1][15:0]),
				 .hw_cos_val_16_1_V_ap_vld(),
				 .hw_cos_val_16_2_V(hw_cos_val_16[2][15:0]),
				 .hw_cos_val_16_2_V_ap_vld(),
				 .hw_cos_val_16_3_V(hw_cos_val_16[3][15:0]),
				 .hw_cos_val_16_3_V_ap_vld(),
				 .hw_cos_val_16_4_V(hw_cos_val_16[4][15:0]),
				 .hw_cos_val_16_4_V_ap_vld(),
				 .hw_cos_val_16_5_V(hw_cos_val_16[5][15:0]),
				 .hw_cos_val_16_5_V_ap_vld(),
				 .hw_cos_val_16_6_V(hw_cos_val_16[6][15:0]),
				 .hw_cos_val_16_6_V_ap_vld(),
				 .hw_cos_val_16_7_V(hw_cos_val_16[7][15:0]),
				 .hw_cos_val_16_7_V_ap_vld(),
				 .hw_cos_val_16_8_V(hw_cos_val_16[8][15:0]),
				 .hw_cos_val_16_8_V_ap_vld(),
				 .hw_cos_val_16_9_V(hw_cos_val_16[9][15:0]),
				 .hw_cos_val_16_9_V_ap_vld(),
				 .hw_cos_val_16_10_V(hw_cos_val_16[10][15:0]),
				 .hw_cos_val_16_10_V_ap_vld(),
				 .hw_cos_val_16_11_V(hw_cos_val_16[11][15:0]),
				 .hw_cos_val_16_11_V_ap_vld(),
				 .hw_cos_val_16_12_V(hw_cos_val_16[12][15:0]),
				 .hw_cos_val_16_12_V_ap_vld(),
				 .hw_cos_val_16_13_V(hw_cos_val_16[13][15:0]),
				 .hw_cos_val_16_13_V_ap_vld(),
				 .hw_cos_val_16_14_V(hw_cos_val_16[14][15:0]),
				 .hw_cos_val_16_14_V_ap_vld(),
				 .hw_cos_val_16_15_V(hw_cos_val_16[15][15:0]),
				 .hw_cos_val_16_15_V_ap_vld(),
				 .cos_rom_sel_0_V(cos_rom_sel_reg[0]),
				 .cos_rom_sel_1_V(cos_rom_sel_reg[1]),
				 .cos_rom_sel_2_V(cos_rom_sel_reg[2]),
				 .cos_rom_sel_3_V(cos_rom_sel_reg[3]),
				 .cos_rom_sel_4_V(cos_rom_sel_reg[4]),
				 .cos_rom_sel_5_V(cos_rom_sel_reg[5]),
				 .cos_rom_sel_6_V(cos_rom_sel_reg[6]),
				 .cos_rom_sel_7_V(cos_rom_sel_reg[7]),
				 .cos_rom_sel_8_V(cos_rom_sel_reg[8]),
				 .cos_rom_sel_9_V(cos_rom_sel_reg[9]),
				 .cos_rom_sel_10_V(cos_rom_sel_reg[10]),
				 .cos_rom_sel_11_V(cos_rom_sel_reg[11]),
				 .cos_rom_sel_12_V(cos_rom_sel_reg[12]),
				 .cos_rom_sel_13_V(cos_rom_sel_reg[13]),
				 .cos_rom_sel_14_V(cos_rom_sel_reg[14]),
				 .cos_rom_sel_15_V(cos_rom_sel_reg[15])
				 );
