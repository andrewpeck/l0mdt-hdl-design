psundara@uciatlaslab.ps.uci.edu.12978:1674253422