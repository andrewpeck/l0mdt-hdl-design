library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;

package l0mdt_dataformats_pkg is

end package l0mdt_dataformats_pkg;

------------------------------------------------------------

package body l0mdt_dataformats_pkg is

end package body l0mdt_dataformats_pkg;
