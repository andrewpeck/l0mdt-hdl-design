psundara@uclhc-2.ps.uci.edu.1286343:1667600067