ilongari@uciatlaslab.ps.uci.edu.31667:1683913032