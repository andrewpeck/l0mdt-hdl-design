--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Guillermo Loustau de Linares             
--  guillermo.ldl@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: drift_time to radius calculation 
--  Description: Autogenerated file          
--     Original File: ../RTInputs/rtdata/rt_pub_run01678_cycle0004_20090422_190058.dat
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package mdt_dt2r_large is

  constant DT2R_LARGE_ADDR_LEN : integer := 10;
  -- constant DT2R_LARGE_DATA_LEN : integer := 9;
  constant DT2R_LARGE_MEM_SIZE : integer := 1024;

  type dt2r_mem_array is array (0 to DT2R_LARGE_MEM_SIZE-1) of integer;
  constant dt2r_large_data : dt2r_mem_array := (
    0 to 8 =>9,
    9 to 18 =>14,
    19 to 28 =>24,
    29 to 38 =>35,
    39 to 48 =>47,
    49 to 58 =>59,
    59 to 68 =>71,
    69 to 78 =>83,
    79 to 88 =>95,
    89 to 98 =>107,
    99 to 108 =>118,
    109 to 118 =>129,
    119 to 128 =>139,
    129 to 138 =>148,
    139 to 148 =>157,
    149 to 158 =>166,
    159 to 168 =>173,
    169 to 178 =>181,
    179 to 188 =>188,
    189 to 198 =>195,
    199 to 208 =>201,
    209 to 218 =>208,
    219 to 228 =>214,
    229 to 238 =>220,
    239 to 248 =>225,
    249 to 258 =>231,
    259 to 268 =>236,
    269 to 278 =>241,
    279 to 288 =>246,
    289 to 298 =>251,
    299 to 308 =>256,
    309 to 318 =>261,
    319 to 328 =>265,
    329 to 338 =>270,
    339 to 348 =>274,
    349 to 358 =>278,
    359 to 368 =>283,
    369 to 378 =>287,
    379 to 388 =>291,
    389 to 398 =>295,
    399 to 408 =>299,
    409 to 418 =>303,
    419 to 428 =>306,
    429 to 438 =>310,
    439 to 448 =>314,
    449 to 458 =>317,
    459 to 468 =>321,
    469 to 477 =>324,
    478 to 487 =>328,
    488 to 497 =>331,
    498 to 507 =>335,
    508 to 517 =>338,
    518 to 527 =>341,
    528 to 537 =>345,
    538 to 547 =>348,
    548 to 557 =>351,
    558 to 567 =>354,
    568 to 577 =>357,
    578 to 587 =>360,
    588 to 597 =>363,
    598 to 607 =>366,
    608 to 617 =>369,
    618 to 627 =>372,
    628 to 637 =>375,
    638 to 647 =>378,
    648 to 657 =>381,
    658 to 667 =>384,
    668 to 677 =>387,
    678 to 687 =>390,
    688 to 697 =>392,
    698 to 707 =>395,
    708 to 717 =>398,
    718 to 727 =>401,
    728 to 737 =>403,
    738 to 747 =>406,
    748 to 757 =>409,
    758 to 767 =>411,
    768 to 777 =>414,
    778 to 787 =>416,
    788 to 797 =>419,
    798 to 807 =>422,
    808 to 817 =>424,
    818 to 827 =>427,
    828 to 837 =>429,
    838 to 847 =>432,
    848 to 857 =>434,
    858 to 867 =>437,
    868 to 877 =>439,
    878 to 887 =>441,
    888 to 897 =>444,
    898 to 907 =>446,
    908 to 917 =>449,
    918 to 927 =>451,
    928 to 937 =>453,
    938 to 946 =>455,
    947 to 956 =>457,
    957 to 966 =>459,
    967 to 976 =>462,
    977 to 1023 =>464 -- original was 987 but simulation gives numbers higher than 987 with very low rate, so we are in hte limit
                      -- I saturate 987 to 1023 until we do more precioson calculations
  );

 end package mdt_dt2r_large;
