--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: rpc_z to tube windows 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package RoI_LUT_BMLA3 is

    type trLUT_limits_t is array (0 to 1) of integer;
    
    type trLUT_layer_t is array (0 to 5) of trLUT_limits_t; -- 1 layer has up to 305 z position
    
    type trLUT_station_t is array (0 to 9130) of trLUT_layer_t; -- 1 station has up to 6 layers

    -- type trLut_sector_t is array ( 0 to 3) of trLUT_station_t; -- 1 sector has 4 station

    constant trLUT_s3m_rom_mem : trLUT_station_t := (
      0 to 30 => ((-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1),(-1,-1)),  
      30 to 60 => ((0,0),(0,0),(0,0),(0,1),(0,1),(0,1)),  
      60 to 90 => ((0,1),(0,1),(0,1),(0,2),(0,2),(0,2)),  
      90 to 120 => ((0,2),(0,2),(0,2),(0,3),(0,3),(0,3)),  
      120 to 150 => ((0,3),(0,3),(0,3),(0,4),(0,4),(0,4)),  
      150 to 180 => ((0,4),(0,4),(0,4),(0,5),(0,5),(0,5)),  
      180 to 210 => ((0,5),(0,5),(0,5),(0,6),(0,6),(0,6)),  
      210 to 240 => ((0,6),(0,6),(0,6),(0,7),(0,7),(0,7)),  
      240 to 270 => ((0,7),(0,7),(0,7),(0,8),(0,8),(0,8)),  
      270 to 300 => ((0,8),(0,8),(0,8),(0,9),(0,9),(0,9)),  
      300 to 330 => ((0,9),(0,9),(0,9),(0,10),(0,10),(0,10)),  
      330 to 360 => ((0,10),(0,10),(0,10),(1,11),(1,11),(1,11)),  
      360 to 390 => ((1,11),(1,11),(1,11),(2,12),(2,12),(2,12)),  
      390 to 420 => ((2,12),(2,12),(2,12),(3,13),(3,13),(3,13)),  
      420 to 450 => ((3,13),(3,13),(3,13),(4,14),(4,14),(4,14)),  
      450 to 480 => ((4,14),(4,14),(4,14),(5,15),(5,15),(5,15)),  
      480 to 510 => ((5,15),(5,15),(5,15),(6,16),(6,16),(6,16)),  
      510 to 540 => ((6,16),(6,16),(6,16),(7,17),(7,17),(7,17)),  
      540 to 570 => ((7,17),(7,17),(7,17),(8,18),(8,18),(9,19)),  
      570 to 600 => ((7,17),(8,18),(8,18),(9,19),(9,19),(10,20)),  
      600 to 630 => ((8,18),(8,18),(9,19),(10,20),(11,21),(11,21)),  
      630 to 660 => ((9,19),(9,19),(10,20),(11,21),(12,22),(12,22)),  
      660 to 690 => ((10,20),(10,20),(10,20),(13,23),(13,23),(13,23)),  
      690 to 720 => ((11,21),(11,21),(11,21),(14,24),(14,24),(14,24)),  
      720 to 750 => ((12,22),(12,22),(12,22),(15,25),(15,25),(15,25)),  
      750 to 780 => ((13,23),(13,23),(13,23),(16,26),(16,26),(16,26)),  
      780 to 810 => ((14,24),(14,24),(14,24),(17,27),(17,27),(17,27)),  
      810 to 840 => ((15,25),(15,25),(15,25),(18,28),(18,28),(18,28)),  
      840 to 870 => ((16,26),(16,26),(16,26),(19,29),(19,29),(19,29)),  
      870 to 900 => ((17,27),(17,27),(17,27),(20,30),(20,30),(20,30)),  
      900 to 930 => ((18,28),(18,28),(18,28),(21,31),(21,31),(21,31)),  
      930 to 960 => ((19,29),(19,29),(19,29),(22,32),(22,32),(22,32)),  
      960 to 990 => ((20,30),(20,30),(20,30),(23,33),(23,33),(23,33)),  
      990 to 1020 => ((21,31),(21,31),(21,31),(24,34),(24,34),(24,34)),  
      1020 to 1050 => ((22,32),(22,32),(22,32),(25,35),(25,35),(25,35)),  
      1050 to 1080 => ((23,33),(23,33),(23,33),(26,36),(26,36),(26,36)),  
      1080 to 1110 => ((24,34),(24,34),(24,34),(27,37),(27,37),(28,38)),  
      1110 to 1140 => ((24,34),(25,35),(25,35),(28,38),(28,38),(29,39)),  
      1140 to 1170 => ((25,35),(26,36),(26,36),(29,39),(29,39),(30,40)),  
      1170 to 1200 => ((26,36),(27,37),(27,37),(30,40),(31,41),(31,41)),  
      1200 to 1230 => ((27,37),(28,38),(28,38),(31,41),(32,42),(32,42)),  
      1230 to 1260 => ((28,38),(28,38),(29,39),(32,42),(33,43),(33,43)),  
      1260 to 1290 => ((29,39),(29,39),(30,40),(33,43),(34,44),(34,44)),  
      1290 to 1320 => ((30,40),(30,40),(31,41),(35,45),(35,45),(35,45)),  
      1320 to 1350 => ((31,41),(31,41),(31,41),(36,46),(36,46),(36,46)),  
      1350 to 1380 => ((32,42),(32,42),(32,42),(37,47),(37,47),(37,47)),  
      1380 to 1410 => ((33,43),(33,43),(33,43),(38,48),(38,48),(38,48)),  
      1410 to 1440 => ((34,44),(34,44),(34,44),(39,49),(39,49),(39,49)),  
      1440 to 1470 => ((35,45),(35,45),(35,45),(40,50),(40,50),(40,50)),  
      1470 to 1500 => ((36,46),(36,46),(36,46),(41,51),(41,51),(41,51)),  
      1500 to 1530 => ((37,47),(37,47),(37,47),(42,52),(42,52),(42,52)),  
      1530 to 1560 => ((38,48),(38,48),(38,48),(43,53),(43,53),(43,53)),  
      1560 to 1590 => ((39,49),(39,49),(39,49),(44,54),(44,54),(44,54)),  
      1590 to 1620 => ((40,50),(40,50),(40,50),(45,55),(45,55),(45,55)),  
      1620 to 1650 => ((41,51),(41,51),(41,51),(46,56),(46,56),(47,56)),  
      1650 to 1680 => ((42,52),(42,52),(42,52),(47,56),(47,57),(48,57)),  
      1680 to 1710 => ((42,52),(43,53),(43,53),(48,57),(48,58),(49,58)),  
      1710 to 1740 => ((43,53),(44,54),(44,54),(49,58),(49,59),(50,59)),  
      1740 to 1770 => ((44,54),(45,55),(45,55),(50,60),(50,60),(51,60)),  
      1770 to 1800 => ((45,55),(46,56),(46,56),(51,61),(52,61),(52,61)),  
      1800 to 1830 => ((46,56),(47,56),(47,56),(52,62),(53,62),(53,62)),  
      1830 to 1860 => ((47,56),(47,57),(48,57),(53,63),(54,63),(54,63)),  
      1860 to 1890 => ((48,57),(48,58),(49,58),(54,64),(55,64),(55,64)),  
      1890 to 1920 => ((49,58),(49,59),(50,59),(55,65),(56,65),(56,65)),  
      1920 to 1950 => ((50,59),(50,60),(51,60),(56,66),(56,66),(56,66)),  
      1950 to 1980 => ((51,60),(51,61),(52,61),(57,67),(57,67),(57,67)),  
      1980 to 2010 => ((52,61),(52,61),(52,62),(58,68),(58,68),(58,68)),  
      2010 to 2040 => ((53,62),(53,62),(53,63),(59,69),(59,69),(60,70)),  
      2040 to 2070 => ((54,63),(54,63),(54,64),(60,70),(60,70),(61,71)),  
      2070 to 2100 => ((55,64),(55,64),(55,65),(61,71),(61,71),(62,72)),  
      2100 to 2130 => ((56,65),(56,65),(56,66),(62,72),(62,72),(63,73)),  
      2130 to 2160 => ((56,66),(56,66),(57,67),(63,73),(63,73),(64,74)),  
      2160 to 2190 => ((57,67),(57,67),(57,67),(64,74),(64,74),(65,75)),  
      2190 to 2220 => ((58,68),(58,68),(58,68),(65,75),(66,76),(66,76)),  
      2220 to 2250 => ((59,69),(59,69),(59,69),(66,76),(67,77),(67,77)),  
      2250 to 2280 => ((60,70),(60,70),(60,70),(67,77),(68,78),(68,78)),  
      2280 to 2310 => ((61,71),(61,71),(61,71),(68,78),(69,79),(69,79)),  
      2310 to 2340 => ((62,72),(62,72),(62,72),(69,79),(70,80),(70,80)),  
      2340 to 2370 => ((63,73),(63,73),(63,73),(70,80),(71,81),(71,81)),  
      2370 to 2400 => ((64,74),(64,74),(64,74),(72,82),(72,82),(72,82)),  
      2400 to 2430 => ((64,74),(65,75),(65,75),(73,83),(73,83),(73,83)),  
      2430 to 2460 => ((65,75),(66,76),(66,76),(74,84),(74,84),(74,84)),  
      2460 to 2490 => ((66,76),(67,77),(67,77),(75,85),(75,85),(75,85)),  
      2490 to 2520 => ((67,77),(68,78),(68,78),(76,86),(76,86),(76,86)),  
      2520 to 2550 => ((68,78),(69,79),(69,79),(77,87),(77,87),(77,87)),  
      2550 to 2580 => ((69,79),(70,80),(70,80),(78,88),(78,88),(79,89)),  
      2580 to 2610 => ((70,80),(70,80),(71,81),(79,89),(79,89),(80,90)),  
      2610 to 2640 => ((71,81),(71,81),(72,82),(80,90),(80,90),(81,91)),  
      2640 to 2670 => ((72,82),(72,82),(73,83),(81,91),(81,91),(82,92)),  
      2670 to 2700 => ((73,83),(73,83),(74,84),(82,92),(82,92),(83,93)),  
      2700 to 2730 => ((74,84),(74,84),(75,85),(83,93),(83,93),(84,94)),  
      2730 to 2760 => ((75,85),(75,85),(76,86),(84,94),(84,94),(85,95)),  
      2760 to 2790 => ((76,86),(76,86),(77,87),(85,95),(86,96),(86,96)),  
      2790 to 2820 => ((77,87),(77,87),(78,88),(86,96),(87,97),(87,97)),  
      2820 to 2850 => ((78,88),(78,88),(78,88),(87,97),(88,98),(88,98)),  
      2850 to 2880 => ((79,89),(79,89),(79,89),(88,98),(89,99),(89,99)),  
      2880 to 2910 => ((80,90),(80,90),(80,90),(89,99),(90,100),(90,100)),  
      2910 to 2940 => ((81,91),(81,91),(81,91),(90,100),(91,101),(91,101)),  
      2940 to 2970 => ((81,91),(82,92),(82,92),(91,101),(92,102),(92,102)),  
      2970 to 3000 => ((82,92),(83,93),(83,93),(92,102),(93,103),(93,103)),  
      3000 to 3030 => ((83,93),(84,94),(84,94),(94,104),(94,104),(94,104)),  
      3030 to 3060 => ((84,94),(85,95),(85,95),(95,105),(95,105),(95,105)),  
      3060 to 3090 => ((85,95),(86,96),(86,96),(96,106),(96,106),(96,106)),  
      3090 to 3120 => ((86,96),(87,97),(87,97),(97,107),(97,107),(98,108)),  
      3120 to 3150 => ((87,97),(88,98),(88,98),(98,108),(98,108),(99,109)),  
      3150 to 3180 => ((88,98),(89,99),(89,99),(99,109),(99,109),(100,110)),  
      3180 to 3210 => ((89,99),(89,99),(90,100),(100,110),(100,110),(101,111)),  
      3210 to 3240 => ((90,100),(90,100),(91,101),(101,111),(101,111),(102,112)),  
      3240 to 3270 => ((91,101),(91,101),(92,102),(102,112),(102,112),(103,112)),  
      3270 to 3300 => ((92,102),(92,102),(93,103),(103,112),(103,113),(104,113)),  
      3300 to 3330 => ((93,103),(93,103),(94,104),(104,113),(104,114),(105,114)),  
      3330 to 3360 => ((94,104),(94,104),(95,105),(105,114),(106,115),(106,115)),  
      3360 to 3390 => ((95,105),(95,105),(96,106),(106,115),(107,116),(107,116)),  
      3390 to 3420 => ((96,106),(96,106),(97,107),(107,116),(108,117),(108,117)),  
      3420 to 3450 => ((97,107),(97,107),(98,108),(108,117),(109,118),(109,118)),  
      3450 to 3480 => ((98,108),(98,108),(99,109),(109,119),(110,119),(110,119)),  
      3480 to 3510 => ((99,109),(99,109),(99,109),(110,120),(111,120),(111,121)),  
      3510 to 3540 => ((99,109),(100,110),(100,110),(111,121),(112,121),(112,122)),  
      3540 to 3570 => ((100,110),(101,111),(101,111),(112,122),(112,122),(113,123)),  
      3570 to 3600 => ((101,111),(102,112),(102,112),(113,123),(113,123),(114,124)),  
      3600 to 3630 => ((102,112),(103,112),(103,113),(114,124),(114,124),(115,125)),  
      3630 to 3660 => ((103,113),(104,113),(104,114),(115,125),(115,125),(116,126)),  
      3660 to 3690 => ((104,113),(105,114),(105,114),(116,126),(116,126),(117,127)),  
      3690 to 3720 => ((105,114),(106,115),(106,115),(117,127),(117,127),(118,128)),  
      3720 to 3750 => ((106,115),(107,116),(107,116),(118,128),(118,128),(119,129)),  
      3750 to 3780 => ((107,116),(108,117),(108,117),(119,129),(120,130),(120,130)),  
      3780 to 3810 => ((108,117),(109,118),(109,118),(120,130),(121,131),(121,131)),  
      3810 to 3840 => ((109,118),(109,119),(110,119),(121,131),(122,132),(122,132)),  
      3840 to 3870 => ((110,119),(110,120),(111,120),(122,132),(123,133),(123,133)),  
      3870 to 3900 => ((111,120),(111,121),(112,121),(123,133),(124,134),(124,134)),  
      3900 to 3930 => ((112,121),(112,122),(112,122),(124,134),(125,135),(125,135)),  
      3930 to 3960 => ((112,122),(113,123),(113,123),(125,135),(126,136),(126,136)),  
      3960 to 3990 => ((113,123),(113,123),(114,124),(126,136),(127,137),(127,137)),  
      3990 to 4020 => ((114,124),(114,124),(115,125),(127,137),(128,138),(128,138)),  
      4020 to 4050 => ((115,125),(115,125),(116,126),(128,138),(129,139),(130,140)),  
      4050 to 4080 => ((116,126),(116,126),(117,127),(129,139),(130,140),(131,141)),  
      4080 to 4110 => ((117,127),(117,127),(118,128),(131,141),(131,141),(132,142)),  
      4110 to 4140 => ((118,128),(118,128),(119,129),(132,142),(132,142),(133,143)),  
      4140 to 4170 => ((119,129),(119,129),(120,130),(133,143),(133,143),(134,144)),  
      4170 to 4200 => ((120,130),(120,130),(121,131),(134,144),(134,144),(135,145)),  
      4200 to 4230 => ((120,130),(121,131),(122,132),(135,145),(135,145),(136,146)),  
      4230 to 4260 => ((121,131),(122,132),(123,133),(136,146),(136,146),(137,147)),  
      4260 to 4290 => ((122,132),(123,133),(124,134),(137,147),(137,147),(138,148)),  
      4290 to 4320 => ((123,133),(124,134),(125,135),(138,148),(138,148),(139,149)),  
      4320 to 4350 => ((124,134),(125,135),(125,135),(139,149),(140,150),(140,150)),  
      4350 to 4380 => ((125,135),(126,136),(126,136),(140,150),(141,151),(141,151)),  
      4380 to 4410 => ((126,136),(127,137),(127,137),(141,151),(142,152),(142,152)),  
      4410 to 4440 => ((127,137),(128,138),(128,138),(142,152),(143,153),(143,153)),  
      4440 to 4470 => ((128,138),(129,139),(129,139),(143,153),(144,154),(144,154)),  
      4470 to 4500 => ((129,139),(130,140),(130,140),(144,154),(145,155),(145,155)),  
      4500 to 4530 => ((130,140),(131,141),(131,141),(145,155),(146,156),(146,156)),  
      4530 to 4560 => ((131,141),(132,142),(132,142),(146,156),(147,157),(147,157)),  
      4560 to 4590 => ((132,142),(132,142),(133,143),(147,157),(148,158),(149,159)),  
      4590 to 4620 => ((133,143),(133,143),(134,144),(148,158),(149,159),(150,160)),  
      4620 to 4650 => ((134,144),(134,144),(135,145),(149,159),(150,160),(151,161)),  
      4650 to 4680 => ((135,145),(135,145),(136,146),(150,160),(151,161),(152,162)),  
      4680 to 4710 => ((136,146),(136,146),(137,147),(151,161),(152,162),(153,163)),  
      4710 to 4740 => ((137,147),(137,147),(138,148),(153,163),(153,163),(154,164)),  
      4740 to 4770 => ((138,148),(138,148),(139,149),(154,164),(154,164),(155,165)),  
      4770 to 4800 => ((138,148),(139,149),(140,150),(155,165),(155,165),(156,166)),  
      4800 to 4830 => ((139,149),(140,150),(141,151),(156,166),(156,166),(157,167)),  
      4830 to 4860 => ((140,150),(141,151),(142,152),(157,167),(157,167),(158,168)),  
      4860 to 4890 => ((141,151),(142,152),(143,153),(158,168),(158,168),(159,168)),  
      4890 to 4920 => ((142,152),(143,153),(144,154),(159,168),(159,169),(160,169)),  
      4920 to 4950 => ((143,153),(144,154),(145,155),(160,169),(161,170),(161,171)),  
      4950 to 4980 => ((144,154),(145,155),(146,156),(161,170),(162,171),(162,172)),  
      4980 to 5010 => ((145,155),(146,156),(146,156),(162,171),(163,172),(163,173)),  
      5010 to 5040 => ((146,156),(147,157),(147,157),(163,172),(164,173),(164,174)),  
      5040 to 5070 => ((147,157),(148,158),(148,158),(164,173),(165,174),(165,175)),  
      5070 to 5100 => ((148,158),(149,159),(149,159),(165,174),(166,175),(167,176)),  
      5100 to 5130 => ((149,159),(150,160),(150,160),(166,175),(167,176),(168,177)),  
      5130 to 5160 => ((150,160),(151,161),(151,161),(167,176),(168,177),(168,178)),  
      5160 to 5190 => ((151,161),(151,161),(152,162),(168,178),(168,178),(169,179)),  
      5190 to 5220 => ((152,162),(152,162),(153,163),(169,179),(169,179),(170,180)),  
      5220 to 5250 => ((153,163),(153,163),(154,164),(170,180),(170,180),(171,181)),  
      5250 to 5280 => ((154,164),(154,164),(155,165),(171,181),(171,181),(172,182)),  
      5280 to 5310 => ((155,165),(155,165),(156,166),(172,182),(172,182),(173,183)),  
      5310 to 5340 => ((155,165),(156,166),(157,167),(173,183),(173,183),(174,184)),  
      5340 to 5370 => ((156,166),(157,167),(158,168),(174,184),(175,185),(175,185)),  
      5370 to 5400 => ((157,167),(158,168),(159,168),(175,185),(176,186),(176,186)),  
      5400 to 5430 => ((158,168),(159,168),(160,169),(176,186),(177,187),(177,187)),  
      5430 to 5460 => ((159,169),(160,169),(161,170),(177,187),(178,188),(178,188)),  
      5460 to 5490 => ((160,170),(161,170),(162,171),(178,188),(179,189),(180,190)),  
      5490 to 5520 => ((161,170),(162,171),(163,172),(179,189),(180,190),(181,191)),  
      5520 to 5550 => ((162,171),(163,172),(164,173),(180,190),(181,191),(182,192)),  
      5550 to 5580 => ((163,172),(164,173),(165,174),(181,191),(182,192),(183,193)),  
      5580 to 5610 => ((164,173),(165,174),(166,175),(182,192),(183,193),(184,194)),  
      5610 to 5640 => ((165,174),(166,175),(167,176),(183,193),(184,194),(185,195)),  
      5640 to 5670 => ((166,175),(167,176),(167,177),(184,194),(185,195),(186,196)),  
      5670 to 5700 => ((167,176),(168,177),(168,178),(185,195),(186,196),(187,197)),  
      5700 to 5730 => ((168,177),(168,178),(169,179),(186,196),(187,197),(188,198)),  
      5730 to 5760 => ((168,178),(169,179),(170,180),(187,197),(188,198),(189,199)),  
      5760 to 5790 => ((169,179),(170,180),(171,181),(188,198),(189,199),(190,200)),  
      5790 to 5820 => ((170,180),(171,181),(172,182),(190,200),(190,200),(191,201)),  
      5820 to 5850 => ((171,181),(172,182),(172,182),(191,201),(191,201),(192,202)),  
      5850 to 5880 => ((172,182),(173,183),(173,183),(192,202),(192,202),(193,203)),  
      5880 to 5910 => ((173,183),(174,184),(174,184),(193,203),(193,203),(194,204)),  
      5910 to 5940 => ((174,184),(175,185),(175,185),(194,204),(195,205),(195,205)),  
      5940 to 5970 => ((175,185),(175,185),(176,186),(195,205),(196,206),(196,206)),  
      5970 to 6000 => ((176,186),(176,186),(177,187),(196,206),(197,207),(197,207)),  
      6000 to 6030 => ((177,187),(177,187),(178,188),(197,207),(198,208),(199,208)),  
      6030 to 6060 => ((177,187),(178,188),(179,189),(198,208),(199,208),(200,209)),  
      6060 to 6090 => ((178,188),(179,189),(180,190),(199,208),(200,209),(201,210)),  
      6090 to 6120 => ((179,189),(180,190),(181,191),(200,209),(201,210),(202,211)),  
      6120 to 6150 => ((180,190),(181,191),(182,192),(201,210),(202,211),(203,212)),  
      6150 to 6180 => ((181,191),(182,192),(183,193),(202,211),(203,212),(204,213)),  
      6180 to 6210 => ((182,192),(183,193),(184,194),(203,212),(204,213),(205,214)),  
      6210 to 6240 => ((183,193),(184,194),(185,195),(204,213),(205,214),(206,215)),  
      6240 to 6270 => ((184,194),(185,195),(186,196),(205,215),(206,215),(207,216)),  
      6270 to 6300 => ((185,195),(186,196),(187,197),(206,216),(207,216),(208,217)),  
      6300 to 6330 => ((186,196),(187,197),(188,198),(207,217),(208,217),(208,218)),  
      6330 to 6360 => ((187,197),(188,198),(189,199),(208,218),(209,219),(209,219)),  
      6360 to 6390 => ((188,198),(189,199),(190,200),(209,219),(210,220),(210,220)),  
      6390 to 6420 => ((189,199),(190,200),(191,201),(210,220),(211,221),(212,222)),  
      6420 to 6450 => ((190,200),(191,201),(192,202),(211,221),(212,222),(213,223)),  
      6450 to 6480 => ((191,201),(192,202),(193,203),(212,222),(213,223),(214,224)),  
      6480 to 6510 => ((192,202),(193,203),(193,203),(213,223),(214,224),(215,225)),  
      6510 to 6540 => ((193,203),(194,204),(194,204),(214,224),(215,225),(216,226)),  
      6540 to 6570 => ((194,204),(194,204),(195,205),(215,225),(216,226),(217,227)),  
      6570 to 6600 => ((195,205),(195,205),(196,206),(216,226),(217,227),(218,228)),  
      6600 to 6630 => ((195,205),(196,206),(197,207),(217,227),(218,228),(219,229)),  
      6630 to 6660 => ((196,206),(197,207),(198,208),(218,228),(219,229),(220,230)),  
      6660 to 6690 => ((197,207),(198,208),(199,209),(219,229),(220,230),(221,231)),  
      6690 to 6720 => ((198,208),(199,209),(200,209),(220,230),(221,231),(222,232)),  
      6720 to 6750 => ((199,209),(200,209),(201,210),(221,231),(222,232),(223,233)),  
      6750 to 6780 => ((200,209),(201,210),(202,211),(222,232),(223,233),(224,234)),  
      6780 to 6810 => ((201,210),(202,211),(203,212),(223,233),(224,234),(225,235)),  
      6810 to 6840 => ((202,211),(203,212),(204,213),(224,234),(225,235),(226,236)),  
      6840 to 6870 => ((203,212),(204,213),(205,214),(225,235),(226,236),(227,237)),  
      6870 to 6900 => ((204,213),(205,214),(206,215),(227,237),(227,237),(228,238)),  
      6900 to 6930 => ((205,214),(206,215),(207,216),(228,238),(229,239),(229,239)),  
      6930 to 6960 => ((206,215),(207,216),(208,217),(229,239),(230,240),(231,241)),  
      6960 to 6990 => ((207,216),(208,217),(208,218),(230,240),(231,241),(232,242)),  
      6990 to 7020 => ((208,217),(208,218),(209,219),(231,241),(232,242),(233,243)),  
      7020 to 7050 => ((208,218),(209,219),(210,220),(232,242),(233,243),(234,244)),  
      7050 to 7080 => ((209,219),(210,220),(211,221),(233,243),(234,244),(235,245)),  
      7080 to 7110 => ((210,220),(211,221),(212,222),(234,244),(235,245),(236,246)),  
      7110 to 7140 => ((211,221),(212,222),(213,223),(235,245),(236,246),(237,247)),  
      7140 to 7170 => ((212,222),(213,223),(214,224),(236,246),(237,247),(238,248)),  
      7170 to 7200 => ((213,223),(214,224),(215,225),(237,247),(238,248),(239,248)),  
      7200 to 7230 => ((214,224),(215,225),(216,226),(238,248),(239,248),(240,249)),  
      7230 to 7260 => ((215,225),(216,226),(217,227),(239,248),(240,249),(241,250)),  
      7260 to 7290 => ((216,226),(217,227),(218,228),(240,249),(241,250),(242,251)),  
      7290 to 7320 => ((217,227),(218,228),(219,229),(241,250),(242,251),(243,253)),  
      7320 to 7350 => ((217,227),(218,228),(220,230),(242,252),(243,253),(244,254)),  
      7350 to 7380 => ((218,228),(219,229),(220,230),(243,253),(244,254),(245,255)),  
      7380 to 7410 => ((219,229),(220,230),(221,231),(244,254),(245,255),(246,256)),  
      7410 to 7440 => ((220,230),(221,231),(222,232),(245,255),(246,256),(247,257)),  
      7440 to 7470 => ((221,231),(222,232),(223,233),(246,256),(247,257),(248,258)),  
      7470 to 7500 => ((222,232),(223,233),(224,234),(247,257),(248,258),(249,259)),  
      7500 to 7530 => ((223,233),(224,234),(225,235),(248,258),(249,259),(250,260)),  
      7530 to 7560 => ((224,234),(225,235),(226,236),(249,259),(250,260),(251,261)),  
      7560 to 7590 => ((225,235),(226,236),(227,237),(250,260),(251,261),(252,262)),  
      7590 to 7620 => ((226,236),(227,237),(228,238),(251,261),(252,262),(253,263)),  
      7620 to 7650 => ((227,237),(228,238),(229,239),(252,262),(253,263),(254,264)),  
      7650 to 7680 => ((228,238),(229,239),(230,240),(253,263),(254,264),(255,265)),  
      7680 to 7710 => ((229,239),(230,240),(231,241),(254,264),(255,265),(256,266)),  
      7710 to 7740 => ((230,240),(231,241),(232,242),(255,265),(256,266),(257,267)),  
      7740 to 7770 => ((231,241),(232,242),(233,243),(256,266),(257,267),(258,268)),  
      7770 to 7800 => ((232,242),(233,243),(234,244),(257,267),(258,268),(259,269)),  
      7800 to 7830 => ((233,243),(234,244),(235,245),(258,268),(259,269),(260,270)),  
      7830 to 7860 => ((234,244),(235,245),(236,246),(259,269),(260,270),(262,272)),  
      7860 to 7890 => ((234,244),(236,246),(237,247),(260,270),(261,271),(263,273)),  
      7890 to 7920 => ((235,245),(237,247),(238,248),(261,271),(263,273),(264,274)),  
      7920 to 7950 => ((236,246),(237,247),(239,248),(262,272),(264,274),(265,275)),  
      7950 to 7980 => ((237,247),(238,248),(240,249),(264,274),(265,275),(266,276)),  
      7980 to 8010 => ((238,248),(239,249),(241,250),(265,275),(266,276),(267,277)),  
      8010 to 8040 => ((239,249),(240,250),(241,251),(266,276),(267,277),(268,278)),  
      8040 to 8070 => ((240,249),(241,251),(242,252),(267,277),(268,278),(269,279)),  
      8070 to 8100 => ((241,250),(242,252),(243,253),(268,278),(269,279),(270,280)),  
      8100 to 8130 => ((242,251),(243,252),(244,254),(269,279),(270,280),(271,281)),  
      8130 to 8160 => ((243,252),(244,253),(245,255),(270,280),(271,281),(272,282)),  
      8160 to 8190 => ((244,253),(245,254),(246,256),(271,281),(272,282),(273,283)),  
      8190 to 8220 => ((245,254),(246,255),(247,256),(272,282),(273,283),(274,284)),  
      8220 to 8250 => ((246,255),(247,256),(248,257),(273,283),(274,284),(275,285)),  
      8250 to 8280 => ((247,256),(248,257),(248,258),(274,284),(275,285),(276,286)),  
      8280 to 8310 => ((248,257),(248,258),(249,259),(275,285),(276,286),(277,287)),  
      8310 to 8340 => ((248,258),(249,259),(250,260),(276,286),(277,287),(278,288)),  
      8340 to 8370 => ((249,259),(250,260),(251,261),(277,287),(278,288),(279,289)),  
      8370 to 8400 => ((250,260),(251,261),(252,262),(278,288),(279,289),(281,291)),  
      8400 to 8430 => ((251,261),(252,262),(253,263),(279,289),(280,290),(282,292)),  
      8430 to 8460 => ((252,262),(253,263),(254,264),(280,290),(281,291),(283,293)),  
      8460 to 8490 => ((253,263),(254,264),(255,265),(281,291),(283,293),(284,294)),  
      8490 to 8520 => ((254,264),(255,265),(256,266),(282,292),(284,294),(285,295)),  
      8520 to 8550 => ((255,265),(256,266),(257,267),(283,293),(285,295),(286,296)),  
      8550 to 8580 => ((256,266),(257,267),(258,268),(284,294),(286,296),(287,297)),  
      8580 to 8610 => ((256,266),(258,268),(259,269),(286,296),(287,297),(288,298)),  
      8610 to 8640 => ((257,267),(259,269),(260,270),(287,297),(288,298),(289,299)),  
      8640 to 8670 => ((258,268),(260,270),(261,271),(288,298),(289,299),(290,300)),  
      8670 to 8700 => ((259,269),(261,271),(262,272),(289,299),(290,300),(291,301)),  
      8700 to 8730 => ((260,270),(261,271),(263,273),(290,300),(291,301),(292,302)),  
      8730 to 8760 => ((261,271),(262,272),(264,274),(291,301),(292,302),(293,303)),  
      8760 to 8790 => ((262,272),(263,273),(265,275),(292,302),(293,303),(294,304)),  
      8790 to 8820 => ((263,273),(264,274),(266,276),(293,303),(294,304),(295,305)),  
      8820 to 8850 => ((264,274),(265,275),(267,277),(294,304),(295,305),(296,306)),  
      8850 to 8880 => ((265,275),(266,276),(267,277),(295,305),(296,306),(297,307)),  
      8880 to 8910 => ((266,276),(267,277),(268,278),(296,306),(297,307),(298,308)),  
      8910 to 8940 => ((267,277),(268,278),(269,279),(297,307),(298,308),(300,310)),  
      8940 to 8970 => ((268,278),(269,279),(270,280),(298,308),(299,309),(301,311)),  
      8970 to 9000 => ((269,279),(270,280),(271,281),(299,309),(300,310),(302,312)),  
      9000 to 9030 => ((270,280),(271,281),(272,282),(300,310),(301,311),(303,313)),  
      9030 to 9060 => ((271,281),(272,282),(273,283),(301,311),(302,312),(304,314)),  
      9060 to 9090 => ((272,282),(273,283),(274,284),(302,312),(304,314),(305,315)),  
      9090 to 9130 => ((273,283),(274,284),(275,285),(303,313),(305,315),(306,316))
  );

 end package RoI_LUT_BMLA3;
