--------------------------------------------------------------------------------
-- Prototype of functions to convert values to/from text for testbenches
--------------------------------------------------------------------------------
-- original   : Eric Hazen
--      v0.1  : GLdL   : added support for TAR
--      v0.2  : GLdL   : moved to ult module

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;
use shared_lib.config_pkg.all;
-- use shared_lib.vhdl2008_functions_pkg.all;
use shared_lib.detector_param_pkg.all;

library ult_lib;
use ult_lib.ult_tb_sim_pkg.all;

package ult_textio_wr_mpl2pt_pkg is

end ult_textio_wr_mpl2pt_pkg;


package body ult_textio_wr_mpl2pt_pkg is

end ult_textio_wr_mpl2pt_pkg;