--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: rpc_z to tube windows 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package RoI_LUT_BOLA3 is

    type trLUT_limits_t is array (0 to 1) of integer;
    
    type trLUT_layer_t is array (0 to 5) of trLUT_limits_t; -- 1 layer has up to 409 z position
    
    type trLUT_station_t is array (0 to 12250) of trLUT_layer_t; -- 1 station has up to 6 layers

    -- type trLut_sector_t is array ( 0 to 3) of trLUT_station_t; -- 1 sector has 4 station

    constant trLUT_s3o_rom_mem : trLUT_station_t := (
      0 to 30 => ((0,1),(0,1),(0,1),(0,1),(0,1),(0,1)),  
      30 to 60 => ((0,2),(0,2),(0,2),(0,3),(0,3),(0,3)),  
      60 to 90 => ((0,3),(0,3),(0,3),(0,4),(0,4),(0,4)),  
      90 to 120 => ((0,4),(0,4),(0,4),(0,5),(0,5),(0,5)),  
      120 to 150 => ((0,5),(0,5),(0,5),(0,6),(0,6),(0,6)),  
      150 to 180 => ((0,6),(0,6),(0,6),(0,7),(0,7),(0,7)),  
      180 to 210 => ((0,7),(0,7),(0,7),(0,8),(0,8),(0,8)),  
      210 to 240 => ((0,8),(0,8),(0,8),(0,9),(0,9),(0,9)),  
      240 to 270 => ((0,9),(0,9),(0,9),(0,10),(0,10),(0,10)),  
      270 to 300 => ((0,10),(0,10),(0,10),(0,11),(0,11),(0,11)),  
      300 to 330 => ((0,11),(0,11),(0,11),(0,12),(0,12),(0,12)),  
      330 to 360 => ((0,12),(0,12),(0,12),(0,13),(0,13),(0,13)),  
      360 to 390 => ((0,13),(0,13),(0,13),(0,14),(0,14),(0,14)),  
      390 to 420 => ((0,14),(0,14),(0,14),(1,15),(1,15),(1,15)),  
      420 to 450 => ((1,15),(1,15),(1,15),(2,16),(2,16),(2,16)),  
      450 to 480 => ((2,16),(2,16),(2,16),(3,17),(3,17),(3,17)),  
      480 to 510 => ((3,17),(3,17),(3,17),(4,18),(4,18),(4,18)),  
      510 to 540 => ((4,18),(4,18),(4,18),(5,19),(5,19),(5,19)),  
      540 to 570 => ((5,19),(5,19),(5,19),(6,20),(6,20),(6,20)),  
      570 to 600 => ((6,20),(6,20),(6,20),(7,21),(7,21),(7,21)),  
      600 to 630 => ((7,21),(7,21),(7,21),(8,22),(8,22),(8,22)),  
      630 to 660 => ((8,22),(8,22),(8,22),(9,23),(9,23),(9,23)),  
      660 to 690 => ((9,23),(9,23),(9,23),(10,24),(10,24),(10,24)),  
      690 to 720 => ((10,24),(10,24),(10,24),(11,25),(11,25),(11,25)),  
      720 to 750 => ((11,25),(11,25),(11,25),(12,26),(12,26),(13,27)),  
      750 to 780 => ((11,25),(12,26),(12,26),(13,27),(13,27),(14,28)),  
      780 to 810 => ((12,26),(13,27),(13,27),(14,28),(15,29),(15,29)),  
      810 to 840 => ((13,27),(13,27),(14,28),(15,29),(16,30),(16,30)),  
      840 to 870 => ((14,28),(14,28),(15,29),(17,31),(17,31),(17,31)),  
      870 to 900 => ((15,29),(15,29),(15,29),(18,32),(18,32),(18,32)),  
      900 to 930 => ((16,30),(16,30),(16,30),(19,33),(19,33),(19,33)),  
      930 to 960 => ((17,31),(17,31),(17,31),(20,34),(20,34),(20,34)),  
      960 to 990 => ((18,32),(18,32),(18,32),(21,35),(21,35),(21,35)),  
      990 to 1020 => ((19,33),(19,33),(19,33),(22,36),(22,36),(22,36)),  
      1020 to 1050 => ((20,34),(20,34),(20,34),(23,37),(23,37),(23,37)),  
      1050 to 1080 => ((21,35),(21,35),(21,35),(24,38),(24,38),(24,38)),  
      1080 to 1110 => ((22,36),(22,36),(22,36),(25,39),(25,39),(25,39)),  
      1110 to 1140 => ((23,37),(23,37),(23,37),(26,40),(26,40),(26,40)),  
      1140 to 1170 => ((24,38),(24,38),(24,38),(27,41),(27,41),(27,41)),  
      1170 to 1200 => ((25,39),(25,39),(25,39),(28,42),(28,42),(28,42)),  
      1200 to 1230 => ((26,40),(26,40),(26,40),(29,43),(29,43),(29,43)),  
      1230 to 1260 => ((27,41),(27,41),(27,41),(30,44),(30,44),(30,44)),  
      1260 to 1290 => ((28,42),(28,42),(28,42),(31,45),(31,45),(31,45)),  
      1290 to 1320 => ((29,43),(29,43),(29,43),(32,46),(32,46),(32,46)),  
      1320 to 1350 => ((30,44),(30,44),(30,44),(33,47),(33,47),(33,47)),  
      1350 to 1380 => ((31,45),(31,45),(31,45),(34,48),(34,48),(34,48)),  
      1380 to 1410 => ((32,46),(32,46),(32,46),(35,49),(35,49),(35,49)),  
      1410 to 1440 => ((33,47),(33,47),(33,47),(36,50),(36,50),(37,51)),  
      1440 to 1470 => ((34,48),(34,48),(34,48),(37,51),(37,51),(38,52)),  
      1470 to 1500 => ((34,48),(35,49),(35,49),(38,52),(38,52),(39,53)),  
      1500 to 1530 => ((35,49),(36,50),(36,50),(39,53),(40,54),(40,54)),  
      1530 to 1560 => ((36,50),(37,51),(37,51),(40,54),(41,55),(41,55)),  
      1560 to 1590 => ((37,51),(38,52),(38,52),(41,55),(42,56),(42,56)),  
      1590 to 1620 => ((38,52),(38,52),(39,53),(42,56),(43,57),(43,57)),  
      1620 to 1650 => ((39,53),(39,53),(40,54),(43,57),(44,58),(44,58)),  
      1650 to 1680 => ((40,54),(40,54),(41,55),(45,59),(45,59),(45,59)),  
      1680 to 1710 => ((41,55),(41,55),(42,56),(46,60),(46,60),(46,60)),  
      1710 to 1740 => ((42,56),(42,56),(43,57),(47,61),(47,61),(47,61)),  
      1740 to 1770 => ((43,57),(43,57),(43,57),(48,62),(48,62),(48,62)),  
      1770 to 1800 => ((44,58),(44,58),(44,58),(49,63),(49,63),(49,63)),  
      1800 to 1830 => ((45,59),(45,59),(45,59),(50,64),(50,64),(50,64)),  
      1830 to 1860 => ((46,60),(46,60),(46,60),(51,65),(51,65),(51,65)),  
      1860 to 1890 => ((47,61),(47,61),(47,61),(52,66),(52,66),(52,66)),  
      1890 to 1920 => ((48,62),(48,62),(48,62),(53,67),(53,67),(53,67)),  
      1920 to 1950 => ((49,63),(49,63),(49,63),(54,68),(54,68),(54,68)),  
      1950 to 1980 => ((50,64),(50,64),(50,64),(55,69),(55,69),(55,69)),  
      1980 to 2010 => ((51,65),(51,65),(51,65),(56,70),(56,70),(56,70)),  
      2010 to 2040 => ((52,66),(52,66),(52,66),(57,71),(57,71),(57,71)),  
      2040 to 2070 => ((53,67),(53,67),(53,67),(58,72),(58,72),(58,72)),  
      2070 to 2100 => ((54,68),(54,68),(54,68),(59,72),(59,73),(59,73)),  
      2100 to 2130 => ((55,69),(55,69),(55,69),(60,73),(60,74),(61,74)),  
      2130 to 2160 => ((56,70),(56,70),(56,70),(61,74),(61,75),(62,75)),  
      2160 to 2190 => ((57,71),(57,71),(57,71),(62,75),(62,76),(63,76)),  
      2190 to 2220 => ((57,71),(58,72),(58,72),(63,76),(63,77),(64,77)),  
      2220 to 2250 => ((58,72),(59,72),(59,72),(64,77),(64,78),(65,78)),  
      2250 to 2280 => ((59,73),(60,73),(60,73),(65,79),(66,79),(66,79)),  
      2280 to 2310 => ((60,74),(61,74),(61,74),(66,80),(67,80),(67,80)),  
      2310 to 2340 => ((61,75),(62,75),(62,75),(67,81),(68,81),(68,81)),  
      2340 to 2370 => ((62,76),(63,76),(63,76),(68,82),(69,82),(69,82)),  
      2370 to 2400 => ((63,76),(63,77),(64,77),(69,83),(70,83),(70,83)),  
      2400 to 2430 => ((64,77),(64,78),(65,78),(70,84),(71,84),(71,84)),  
      2430 to 2460 => ((65,78),(65,79),(66,79),(71,85),(72,85),(72,85)),  
      2460 to 2490 => ((66,79),(66,80),(67,80),(72,86),(72,86),(72,86)),  
      2490 to 2520 => ((67,80),(67,81),(68,81),(73,87),(73,87),(73,87)),  
      2520 to 2550 => ((68,81),(68,82),(69,82),(74,88),(74,88),(74,88)),  
      2550 to 2580 => ((69,82),(69,83),(70,83),(75,89),(75,89),(75,89)),  
      2580 to 2610 => ((70,83),(70,83),(70,84),(76,90),(76,90),(76,90)),  
      2610 to 2640 => ((71,84),(71,84),(71,85),(77,91),(77,91),(78,92)),  
      2640 to 2670 => ((72,85),(72,85),(72,86),(78,92),(78,92),(79,93)),  
      2670 to 2700 => ((72,86),(72,86),(73,87),(79,93),(79,93),(80,94)),  
      2700 to 2730 => ((73,87),(73,87),(74,88),(80,94),(80,94),(81,95)),  
      2730 to 2760 => ((74,88),(74,88),(75,89),(81,95),(81,95),(82,96)),  
      2760 to 2790 => ((75,89),(75,89),(76,90),(82,96),(82,96),(83,97)),  
      2790 to 2820 => ((76,90),(76,90),(77,91),(83,97),(83,97),(84,98)),  
      2820 to 2850 => ((77,91),(77,91),(77,91),(84,98),(85,99),(85,99)),  
      2850 to 2880 => ((78,92),(78,92),(78,92),(85,99),(86,100),(86,100)),  
      2880 to 2910 => ((79,93),(79,93),(79,93),(86,100),(87,101),(87,101)),  
      2910 to 2940 => ((80,94),(80,94),(80,94),(87,101),(88,102),(88,102)),  
      2940 to 2970 => ((81,95),(81,95),(81,95),(88,102),(89,103),(89,103)),  
      2970 to 3000 => ((82,96),(82,96),(82,96),(89,103),(90,104),(90,104)),  
      3000 to 3030 => ((83,97),(83,97),(83,97),(90,104),(91,105),(91,105)),  
      3030 to 3060 => ((84,98),(84,98),(84,98),(91,105),(92,106),(92,106)),  
      3060 to 3090 => ((85,99),(85,99),(85,99),(93,107),(93,107),(93,107)),  
      3090 to 3120 => ((85,99),(86,100),(86,100),(94,108),(94,108),(94,108)),  
      3120 to 3150 => ((86,100),(87,101),(87,101),(95,109),(95,109),(95,109)),  
      3150 to 3180 => ((87,101),(88,102),(88,102),(96,110),(96,110),(96,110)),  
      3180 to 3210 => ((88,102),(89,103),(89,103),(97,111),(97,111),(97,111)),  
      3210 to 3240 => ((89,103),(90,104),(90,104),(98,112),(98,112),(98,112)),  
      3240 to 3270 => ((90,104),(91,105),(91,105),(99,113),(99,113),(99,113)),  
      3270 to 3300 => ((91,105),(92,106),(92,106),(100,114),(100,114),(100,114)),  
      3300 to 3330 => ((92,106),(93,107),(93,107),(101,115),(101,115),(102,116)),  
      3330 to 3360 => ((93,107),(94,108),(94,108),(102,116),(102,116),(103,117)),  
      3360 to 3390 => ((94,108),(94,108),(95,109),(103,117),(103,117),(104,118)),  
      3390 to 3420 => ((95,109),(95,109),(96,110),(104,118),(104,118),(105,119)),  
      3420 to 3450 => ((96,110),(96,110),(97,111),(105,119),(105,119),(106,120)),  
      3450 to 3480 => ((97,111),(97,111),(98,112),(106,120),(106,120),(107,121)),  
      3480 to 3510 => ((98,112),(98,112),(99,113),(107,121),(107,121),(108,122)),  
      3510 to 3540 => ((99,113),(99,113),(100,114),(108,122),(108,122),(109,123)),  
      3540 to 3570 => ((100,114),(100,114),(101,115),(109,123),(109,123),(110,124)),  
      3570 to 3600 => ((101,115),(101,115),(102,116),(110,124),(111,125),(111,125)),  
      3600 to 3630 => ((102,116),(102,116),(103,117),(111,125),(112,126),(112,126)),  
      3630 to 3660 => ((103,117),(103,117),(104,118),(112,126),(113,127),(113,127)),  
      3660 to 3690 => ((104,118),(104,118),(104,118),(113,127),(114,128),(114,128)),  
      3690 to 3720 => ((105,119),(105,119),(105,119),(114,128),(115,129),(115,129)),  
      3720 to 3750 => ((106,120),(106,120),(106,120),(115,129),(116,130),(116,130)),  
      3750 to 3780 => ((107,121),(107,121),(107,121),(116,130),(117,131),(117,131)),  
      3780 to 3810 => ((108,122),(108,122),(108,122),(117,131),(118,132),(118,132)),  
      3810 to 3840 => ((109,123),(109,123),(109,123),(118,132),(119,133),(119,133)),  
      3840 to 3870 => ((109,123),(110,124),(110,124),(119,133),(120,134),(120,134)),  
      3870 to 3900 => ((110,124),(111,125),(111,125),(121,135),(121,135),(121,135)),  
      3900 to 3930 => ((111,125),(112,126),(112,126),(122,136),(122,136),(122,136)),  
      3930 to 3960 => ((112,126),(113,127),(113,127),(123,137),(123,137),(123,137)),  
      3960 to 3990 => ((113,127),(114,128),(114,128),(124,138),(124,138),(124,138)),  
      3990 to 4020 => ((114,128),(115,129),(115,129),(125,139),(125,139),(126,140)),  
      4020 to 4050 => ((115,129),(116,130),(116,130),(126,140),(126,140),(127,141)),  
      4050 to 4080 => ((116,130),(117,131),(117,131),(127,141),(127,141),(128,142)),  
      4080 to 4110 => ((117,131),(118,132),(118,132),(128,142),(128,142),(129,143)),  
      4110 to 4140 => ((118,132),(119,133),(119,133),(129,143),(129,143),(130,144)),  
      4140 to 4170 => ((119,133),(119,133),(120,134),(130,144),(130,144),(131,144)),  
      4170 to 4200 => ((120,134),(120,134),(121,135),(131,144),(131,145),(132,145)),  
      4200 to 4230 => ((121,135),(121,135),(122,136),(132,145),(132,146),(133,146)),  
      4230 to 4260 => ((122,136),(122,136),(123,137),(133,146),(133,147),(134,147)),  
      4260 to 4290 => ((123,137),(123,137),(124,138),(134,147),(134,148),(135,148)),  
      4290 to 4320 => ((124,138),(124,138),(125,139),(135,148),(135,149),(136,149)),  
      4320 to 4350 => ((125,139),(125,139),(126,140),(136,149),(137,150),(137,150)),  
      4350 to 4380 => ((126,140),(126,140),(127,141),(137,150),(138,151),(138,151)),  
      4380 to 4410 => ((127,141),(127,141),(128,142),(138,151),(139,152),(139,152)),  
      4410 to 4440 => ((128,142),(128,142),(129,143),(139,152),(140,153),(140,153)),  
      4440 to 4470 => ((129,143),(129,143),(130,144),(140,153),(141,154),(141,154)),  
      4470 to 4500 => ((130,144),(130,144),(131,144),(141,155),(142,155),(142,155)),  
      4500 to 4530 => ((131,144),(131,144),(132,145),(142,156),(143,156),(143,157)),  
      4530 to 4560 => ((132,145),(132,145),(132,146),(143,157),(144,157),(144,158)),  
      4560 to 4590 => ((132,146),(133,146),(133,147),(144,158),(144,158),(145,159)),  
      4590 to 4620 => ((133,147),(134,147),(134,148),(145,159),(145,159),(146,160)),  
      4620 to 4650 => ((134,148),(135,148),(135,149),(146,160),(146,160),(147,161)),  
      4650 to 4680 => ((135,149),(136,149),(136,150),(147,161),(147,161),(148,162)),  
      4680 to 4710 => ((136,150),(137,150),(137,151),(148,162),(148,162),(149,163)),  
      4710 to 4740 => ((137,151),(138,151),(138,152),(149,163),(149,163),(150,164)),  
      4740 to 4770 => ((138,151),(139,152),(139,153),(150,164),(150,164),(151,165)),  
      4770 to 4800 => ((139,152),(140,153),(140,153),(151,165),(151,165),(152,166)),  
      4800 to 4830 => ((140,153),(141,154),(141,154),(152,166),(152,166),(153,167)),  
      4830 to 4860 => ((141,154),(142,155),(142,155),(153,167),(153,167),(154,168)),  
      4860 to 4890 => ((142,155),(143,156),(143,156),(154,168),(155,169),(155,169)),  
      4890 to 4920 => ((143,156),(144,157),(144,157),(155,169),(156,170),(156,170)),  
      4920 to 4950 => ((144,157),(144,158),(144,158),(156,170),(157,171),(157,171)),  
      4950 to 4980 => ((144,158),(145,159),(145,159),(157,171),(158,172),(158,172)),  
      4980 to 5010 => ((145,159),(146,160),(146,160),(158,172),(159,173),(159,173)),  
      5010 to 5040 => ((146,160),(147,161),(147,161),(159,173),(160,174),(160,174)),  
      5040 to 5070 => ((147,161),(148,162),(148,162),(160,174),(161,175),(161,175)),  
      5070 to 5100 => ((148,162),(149,163),(149,163),(161,175),(162,176),(162,176)),  
      5100 to 5130 => ((149,163),(150,164),(150,164),(162,176),(163,177),(163,177)),  
      5130 to 5160 => ((150,164),(150,164),(151,165),(163,177),(164,178),(164,178)),  
      5160 to 5190 => ((151,165),(151,165),(152,166),(164,178),(165,179),(165,179)),  
      5190 to 5220 => ((152,166),(152,166),(153,167),(165,179),(166,180),(167,181)),  
      5220 to 5250 => ((153,167),(153,167),(154,168),(166,180),(167,181),(168,182)),  
      5250 to 5280 => ((154,168),(154,168),(155,169),(167,181),(168,182),(169,183)),  
      5280 to 5310 => ((155,169),(155,169),(156,170),(169,183),(169,183),(170,184)),  
      5310 to 5340 => ((156,170),(156,170),(157,171),(170,184),(170,184),(171,185)),  
      5340 to 5370 => ((157,171),(157,171),(158,172),(171,185),(171,185),(172,186)),  
      5370 to 5400 => ((158,172),(158,172),(159,173),(172,186),(172,186),(173,187)),  
      5400 to 5430 => ((159,173),(159,173),(160,174),(173,187),(173,187),(174,188)),  
      5430 to 5460 => ((160,174),(160,174),(161,175),(174,188),(174,188),(175,189)),  
      5460 to 5490 => ((160,174),(161,175),(162,176),(175,189),(175,189),(176,190)),  
      5490 to 5520 => ((161,175),(162,176),(163,177),(176,190),(176,190),(177,191)),  
      5520 to 5550 => ((162,176),(163,177),(164,178),(177,191),(177,191),(178,192)),  
      5550 to 5580 => ((163,177),(164,178),(165,179),(178,192),(178,192),(179,193)),  
      5580 to 5610 => ((164,178),(165,179),(166,180),(179,193),(179,193),(180,194)),  
      5610 to 5640 => ((165,179),(166,180),(166,180),(180,194),(181,195),(181,195)),  
      5640 to 5670 => ((166,180),(167,181),(167,181),(181,195),(182,196),(182,196)),  
      5670 to 5700 => ((167,181),(168,182),(168,182),(182,196),(183,197),(183,197)),  
      5700 to 5730 => ((168,182),(169,183),(169,183),(183,197),(184,198),(184,198)),  
      5730 to 5760 => ((169,183),(170,184),(170,184),(184,198),(185,199),(185,199)),  
      5760 to 5790 => ((170,184),(171,185),(171,185),(185,199),(186,200),(186,200)),  
      5790 to 5820 => ((171,185),(172,186),(172,186),(186,200),(187,200),(187,201)),  
      5820 to 5850 => ((172,186),(173,187),(173,187),(187,200),(188,201),(188,202)),  
      5850 to 5880 => ((173,187),(174,188),(174,188),(188,201),(189,202),(189,203)),  
      5880 to 5910 => ((174,188),(175,189),(175,189),(189,203),(190,203),(191,204)),  
      5910 to 5940 => ((175,189),(176,190),(176,190),(190,204),(191,204),(192,205)),  
      5940 to 5970 => ((176,190),(176,190),(177,191),(191,205),(192,205),(193,206)),  
      5970 to 6000 => ((177,191),(177,191),(178,192),(192,206),(193,206),(194,207)),  
      6000 to 6030 => ((178,192),(178,192),(179,193),(193,207),(194,207),(195,208)),  
      6030 to 6060 => ((179,193),(179,193),(180,194),(194,208),(195,208),(196,209)),  
      6060 to 6090 => ((180,194),(180,194),(181,195),(195,209),(196,209),(197,210)),  
      6090 to 6120 => ((181,195),(181,195),(182,196),(197,210),(197,210),(198,211)),  
      6120 to 6150 => ((182,196),(182,196),(183,197),(198,211),(198,211),(199,212)),  
      6150 to 6180 => ((183,197),(183,197),(184,198),(199,212),(199,213),(200,213)),  
      6180 to 6210 => ((183,197),(184,198),(185,199),(200,213),(200,214),(200,214)),  
      6210 to 6240 => ((184,198),(185,199),(186,200),(200,214),(201,215),(201,215)),  
      6240 to 6270 => ((185,199),(186,200),(187,200),(201,215),(202,216),(202,216)),  
      6270 to 6300 => ((186,200),(187,200),(188,201),(202,216),(203,217),(203,217)),  
      6300 to 6330 => ((187,201),(188,201),(189,202),(203,217),(204,218),(204,218)),  
      6330 to 6360 => ((188,202),(189,202),(190,203),(204,218),(205,219),(205,219)),  
      6360 to 6390 => ((189,203),(190,203),(191,204),(205,219),(206,220),(206,220)),  
      6390 to 6420 => ((190,203),(191,204),(192,205),(206,220),(207,221),(208,222)),  
      6420 to 6450 => ((191,204),(192,205),(193,206),(207,221),(208,222),(209,223)),  
      6450 to 6480 => ((192,205),(193,206),(194,207),(208,222),(209,223),(210,224)),  
      6480 to 6510 => ((193,206),(194,207),(194,208),(209,223),(210,224),(211,225)),  
      6510 to 6540 => ((194,207),(195,208),(195,209),(210,224),(211,225),(212,226)),  
      6540 to 6570 => ((195,208),(196,209),(196,210),(211,225),(212,226),(213,227)),  
      6570 to 6600 => ((196,209),(197,210),(197,211),(212,226),(213,227),(214,228)),  
      6600 to 6630 => ((197,210),(198,211),(198,212),(213,227),(214,228),(215,229)),  
      6630 to 6660 => ((198,211),(199,212),(199,213),(214,228),(215,229),(216,230)),  
      6660 to 6690 => ((199,212),(200,213),(200,214),(215,229),(216,230),(217,231)),  
      6690 to 6720 => ((200,213),(200,214),(201,215),(217,231),(217,231),(218,232)),  
      6720 to 6750 => ((200,214),(201,215),(201,215),(218,232),(218,232),(219,233)),  
      6750 to 6780 => ((201,215),(202,216),(202,216),(219,233),(219,233),(220,234)),  
      6780 to 6810 => ((202,216),(203,217),(203,217),(220,234),(220,234),(221,235)),  
      6810 to 6840 => ((203,217),(204,218),(204,218),(221,235),(221,235),(222,236)),  
      6840 to 6870 => ((204,218),(205,219),(205,219),(222,236),(222,236),(223,237)),  
      6870 to 6900 => ((205,219),(206,220),(206,220),(223,237),(223,237),(224,238)),  
      6900 to 6930 => ((206,220),(207,221),(207,221),(224,238),(225,239),(225,239)),  
      6930 to 6960 => ((207,221),(207,221),(208,222),(225,239),(226,240),(226,240)),  
      6960 to 6990 => ((208,222),(208,222),(209,223),(226,240),(227,241),(227,241)),  
      6990 to 7020 => ((209,223),(209,223),(210,224),(227,241),(228,242),(228,242)),  
      7020 to 7050 => ((210,224),(210,224),(211,225),(228,242),(229,243),(229,243)),  
      7050 to 7080 => ((211,225),(211,225),(212,226),(229,243),(230,244),(230,244)),  
      7080 to 7110 => ((212,226),(212,226),(213,227),(230,244),(231,245),(232,246)),  
      7110 to 7140 => ((212,226),(213,227),(214,228),(231,245),(232,246),(233,247)),  
      7140 to 7170 => ((213,227),(214,228),(215,229),(232,246),(233,247),(234,248)),  
      7170 to 7200 => ((214,228),(215,229),(216,230),(233,247),(234,248),(235,249)),  
      7200 to 7230 => ((215,229),(216,230),(217,231),(234,248),(235,249),(236,250)),  
      7230 to 7260 => ((216,230),(217,231),(218,232),(235,249),(236,250),(237,251)),  
      7260 to 7290 => ((217,231),(218,232),(219,233),(236,250),(237,251),(238,252)),  
      7290 to 7320 => ((218,232),(219,233),(220,234),(237,251),(238,252),(239,253)),  
      7320 to 7350 => ((219,233),(220,234),(221,235),(238,252),(239,253),(240,254)),  
      7350 to 7380 => ((220,234),(221,235),(222,236),(239,253),(240,254),(241,255)),  
      7380 to 7410 => ((221,235),(222,236),(223,237),(240,254),(241,255),(242,256)),  
      7410 to 7440 => ((222,236),(223,237),(224,238),(241,255),(242,256),(243,257)),  
      7440 to 7470 => ((223,237),(224,238),(225,239),(242,256),(243,257),(244,258)),  
      7470 to 7500 => ((224,238),(225,239),(226,240),(243,257),(244,258),(245,259)),  
      7500 to 7530 => ((225,239),(226,240),(227,241),(245,259),(245,259),(246,260)),  
      7530 to 7560 => ((226,240),(227,241),(228,242),(246,260),(246,260),(247,261)),  
      7560 to 7590 => ((227,241),(228,242),(229,243),(247,261),(247,261),(248,262)),  
      7590 to 7620 => ((228,242),(229,243),(229,243),(248,262),(248,262),(249,263)),  
      7620 to 7650 => ((229,243),(230,244),(230,244),(249,263),(249,263),(250,264)),  
      7650 to 7680 => ((230,244),(231,245),(231,245),(250,264),(251,265),(251,265)),  
      7680 to 7710 => ((231,245),(232,246),(232,246),(251,265),(252,266),(252,266)),  
      7710 to 7740 => ((232,246),(232,246),(233,247),(252,266),(253,267),(253,267)),  
      7740 to 7770 => ((233,247),(233,247),(234,248),(253,267),(254,268),(254,268)),  
      7770 to 7800 => ((234,248),(234,248),(235,249),(254,268),(255,269),(256,270)),  
      7800 to 7830 => ((235,249),(235,249),(236,250),(255,269),(256,270),(257,271)),  
      7830 to 7860 => ((235,249),(236,250),(237,251),(256,270),(257,271),(258,272)),  
      7860 to 7890 => ((236,250),(237,251),(238,252),(257,271),(258,272),(259,272)),  
      7890 to 7920 => ((237,251),(238,252),(239,253),(258,272),(259,272),(260,273)),  
      7920 to 7950 => ((238,252),(239,253),(240,254),(259,272),(260,273),(261,274)),  
      7950 to 7980 => ((239,253),(240,254),(241,255),(260,273),(261,274),(262,275)),  
      7980 to 8010 => ((240,254),(241,255),(242,256),(261,274),(262,275),(263,276)),  
      8010 to 8040 => ((241,255),(242,256),(243,257),(262,275),(263,276),(264,277)),  
      8040 to 8070 => ((242,256),(243,257),(244,258),(263,276),(264,277),(265,278)),  
      8070 to 8100 => ((243,257),(244,258),(245,259),(264,277),(265,278),(266,279)),  
      8100 to 8130 => ((244,258),(245,259),(246,260),(265,279),(266,279),(267,280)),  
      8130 to 8160 => ((245,259),(246,260),(247,261),(266,280),(267,280),(268,281)),  
      8160 to 8190 => ((246,260),(247,261),(248,262),(267,281),(268,281),(269,282)),  
      8190 to 8220 => ((247,261),(248,262),(249,263),(268,282),(269,283),(270,283)),  
      8220 to 8250 => ((248,262),(249,263),(250,264),(269,283),(270,284),(271,284)),  
      8250 to 8280 => ((249,263),(250,264),(251,265),(270,284),(271,285),(272,285)),  
      8280 to 8310 => ((250,264),(251,265),(252,266),(271,285),(272,286),(273,287)),  
      8310 to 8340 => ((251,265),(252,266),(253,267),(272,286),(273,287),(274,288)),  
      8340 to 8370 => ((252,266),(253,267),(254,268),(273,287),(274,288),(275,289)),  
      8370 to 8400 => ((253,267),(254,268),(255,269),(274,288),(275,289),(276,290)),  
      8400 to 8430 => ((254,268),(255,269),(256,270),(275,289),(276,290),(277,291)),  
      8430 to 8460 => ((255,269),(256,270),(256,270),(276,290),(277,291),(278,292)),  
      8460 to 8490 => ((256,270),(257,271),(257,271),(277,291),(278,292),(279,293)),  
      8490 to 8520 => ((257,271),(258,272),(258,272),(278,292),(279,293),(280,294)),  
      8520 to 8550 => ((258,272),(258,272),(259,273),(279,293),(280,294),(281,295)),  
      8550 to 8580 => ((259,272),(259,273),(260,274),(280,294),(281,295),(282,296)),  
      8580 to 8610 => ((259,273),(260,274),(261,275),(281,295),(282,296),(283,297)),  
      8610 to 8640 => ((260,274),(261,275),(262,276),(282,296),(283,297),(284,298)),  
      8640 to 8670 => ((261,275),(262,276),(263,277),(283,297),(284,298),(285,299)),  
      8670 to 8700 => ((262,276),(263,277),(264,277),(284,298),(285,299),(286,300)),  
      8700 to 8730 => ((263,277),(264,277),(265,278),(285,299),(286,300),(287,301)),  
      8730 to 8760 => ((264,278),(265,278),(266,279),(286,300),(287,301),(288,302)),  
      8760 to 8790 => ((265,278),(266,279),(267,280),(287,301),(288,302),(289,303)),  
      8790 to 8820 => ((266,279),(267,280),(268,281),(288,302),(289,303),(290,304)),  
      8820 to 8850 => ((267,280),(268,281),(269,282),(289,303),(290,304),(291,305)),  
      8850 to 8880 => ((268,281),(269,282),(270,283),(290,304),(291,305),(292,306)),  
      8880 to 8910 => ((269,282),(270,283),(271,284),(291,305),(292,306),(293,307)),  
      8910 to 8940 => ((270,283),(271,284),(272,285),(293,307),(293,307),(294,308)),  
      8940 to 8970 => ((271,284),(272,285),(272,286),(294,308),(295,309),(295,309)),  
      8970 to 9000 => ((272,285),(272,286),(273,287),(295,309),(296,310),(297,311)),  
      9000 to 9030 => ((272,286),(273,287),(274,288),(296,310),(297,311),(298,312)),  
      9030 to 9060 => ((273,287),(274,288),(275,289),(297,311),(298,312),(299,313)),  
      9060 to 9090 => ((274,288),(275,289),(276,290),(298,312),(299,313),(300,314)),  
      9090 to 9120 => ((275,289),(276,290),(277,291),(299,313),(300,314),(301,315)),  
      9120 to 9150 => ((276,290),(277,291),(278,292),(300,314),(301,315),(302,316)),  
      9150 to 9180 => ((277,291),(278,292),(279,293),(301,315),(302,316),(303,317)),  
      9180 to 9210 => ((278,292),(279,293),(280,294),(302,316),(303,317),(304,318)),  
      9210 to 9240 => ((279,293),(280,294),(281,295),(303,317),(304,318),(305,319)),  
      9240 to 9270 => ((280,294),(281,295),(282,296),(304,318),(305,319),(306,320)),  
      9270 to 9300 => ((281,295),(282,296),(283,297),(305,319),(306,320),(307,321)),  
      9300 to 9330 => ((282,296),(283,297),(284,298),(306,320),(307,321),(308,322)),  
      9330 to 9360 => ((283,297),(284,298),(285,299),(307,321),(308,322),(309,323)),  
      9360 to 9390 => ((284,298),(285,299),(286,300),(308,322),(309,323),(310,324)),  
      9390 to 9420 => ((285,299),(286,300),(287,301),(309,323),(310,324),(311,325)),  
      9420 to 9450 => ((286,300),(287,301),(288,302),(310,324),(311,325),(312,326)),  
      9450 to 9480 => ((287,301),(288,302),(289,303),(311,325),(312,326),(313,327)),  
      9480 to 9510 => ((287,301),(289,303),(290,304),(312,326),(313,327),(314,328)),  
      9510 to 9540 => ((288,302),(289,303),(290,304),(313,327),(314,328),(315,329)),  
      9540 to 9570 => ((289,303),(290,304),(291,305),(314,328),(315,329),(316,330)),  
      9570 to 9600 => ((290,304),(291,305),(292,306),(315,329),(316,330),(317,331)),  
      9600 to 9630 => ((291,305),(292,306),(293,307),(316,330),(317,331),(318,332)),  
      9630 to 9660 => ((292,306),(293,307),(294,308),(317,331),(318,332),(319,333)),  
      9660 to 9690 => ((293,307),(294,308),(295,309),(318,332),(319,333),(321,335)),  
      9690 to 9720 => ((294,308),(295,309),(296,310),(319,333),(321,335),(322,336)),  
      9720 to 9750 => ((295,309),(296,310),(297,311),(321,335),(322,336),(323,337)),  
      9750 to 9780 => ((296,310),(297,311),(298,312),(322,336),(323,337),(324,338)),  
      9780 to 9810 => ((297,311),(298,312),(299,313),(323,337),(324,338),(325,339)),  
      9810 to 9840 => ((298,312),(299,313),(300,314),(324,338),(325,339),(326,340)),  
      9840 to 9870 => ((299,313),(300,314),(301,315),(325,339),(326,340),(327,341)),  
      9870 to 9900 => ((300,314),(301,315),(302,316),(326,340),(327,341),(328,342)),  
      9900 to 9930 => ((301,315),(302,316),(303,317),(327,341),(328,342),(329,343)),  
      9930 to 9960 => ((302,316),(303,317),(304,318),(328,342),(329,343),(330,344)),  
      9960 to 9990 => ((303,317),(304,318),(305,319),(329,343),(330,344),(331,344)),  
      9990 to 10020 => ((304,318),(305,319),(306,320),(330,344),(331,344),(332,345)),  
      10020 to 10050 => ((305,319),(306,320),(307,321),(331,344),(332,345),(333,346)),  
      10050 to 10080 => ((306,320),(307,321),(308,322),(332,345),(333,346),(334,347)),  
      10080 to 10110 => ((307,321),(308,322),(309,323),(333,346),(334,347),(335,348)),  
      10110 to 10140 => ((308,322),(309,323),(310,324),(334,347),(335,348),(336,349)),  
      10140 to 10170 => ((309,323),(310,324),(311,325),(335,348),(336,349),(337,350)),  
      10170 to 10200 => ((310,324),(311,325),(312,326),(336,349),(337,350),(338,352)),  
      10200 to 10230 => ((310,324),(312,326),(313,327),(337,350),(338,351),(339,353)),  
      10230 to 10260 => ((311,325),(313,327),(314,328),(338,351),(339,352),(340,354)),  
      10260 to 10290 => ((312,326),(314,328),(315,329),(339,352),(340,354),(341,355)),  
      10290 to 10320 => ((313,327),(314,328),(316,330),(340,353),(341,355),(342,356)),  
      10320 to 10350 => ((314,328),(315,329),(317,331),(341,355),(342,356),(343,357)),  
      10350 to 10380 => ((315,329),(316,330),(318,332),(342,356),(343,357),(344,358)),  
      10380 to 10410 => ((316,330),(317,331),(318,332),(343,357),(344,358),(345,359)),  
      10410 to 10440 => ((317,331),(318,332),(319,333),(344,358),(345,359),(346,360)),  
      10440 to 10470 => ((318,332),(319,333),(320,334),(345,359),(346,360),(347,361)),  
      10470 to 10500 => ((319,333),(320,334),(321,335),(346,360),(347,361),(348,362)),  
      10500 to 10530 => ((320,334),(321,335),(322,336),(347,361),(348,362),(349,363)),  
      10530 to 10560 => ((321,335),(322,336),(323,337),(348,362),(349,363),(350,364)),  
      10560 to 10590 => ((322,336),(323,337),(324,338),(349,363),(350,364),(351,365)),  
      10590 to 10620 => ((323,337),(324,338),(325,339),(350,364),(351,365),(352,366)),  
      10620 to 10650 => ((324,338),(325,339),(326,340),(351,365),(352,366),(353,367)),  
      10650 to 10680 => ((325,339),(326,340),(327,341),(352,366),(353,367),(354,368)),  
      10680 to 10710 => ((326,340),(327,341),(328,342),(353,367),(354,368),(355,369)),  
      10710 to 10740 => ((327,341),(328,342),(329,343),(354,368),(355,369),(356,370)),  
      10740 to 10770 => ((328,342),(329,343),(330,344),(355,369),(356,370),(357,371)),  
      10770 to 10800 => ((329,343),(330,344),(331,344),(356,370),(357,371),(358,372)),  
      10800 to 10830 => ((330,344),(331,344),(332,345),(357,371),(358,372),(359,373)),  
      10830 to 10860 => ((331,344),(332,345),(333,346),(358,372),(359,373),(360,374)),  
      10860 to 10890 => ((332,345),(333,346),(334,347),(359,373),(360,374),(362,376)),  
      10890 to 10920 => ((333,346),(334,347),(335,348),(360,374),(361,375),(363,377)),  
      10920 to 10950 => ((333,347),(335,348),(336,349),(361,375),(362,376),(364,378)),  
      10950 to 10980 => ((334,348),(336,349),(337,350),(362,376),(363,377),(365,379)),  
      10980 to 11010 => ((335,349),(337,350),(338,351),(363,377),(365,379),(366,380)),  
      11010 to 11040 => ((336,350),(338,351),(339,352),(364,378),(366,380),(367,381)),  
      11040 to 11070 => ((337,351),(339,352),(340,353),(365,379),(367,381),(368,382)),  
      11070 to 11100 => ((338,352),(339,353),(341,354),(366,380),(368,382),(369,383)),  
      11100 to 11130 => ((339,353),(340,354),(342,355),(367,381),(369,383),(370,384)),  
      11130 to 11160 => ((340,353),(341,355),(343,356),(369,383),(370,384),(371,385)),  
      11160 to 11190 => ((341,354),(342,356),(344,357),(370,384),(371,385),(372,386)),  
      11190 to 11220 => ((342,355),(343,357),(344,358),(371,385),(372,386),(373,387)),  
      11220 to 11250 => ((343,356),(344,358),(345,359),(372,386),(373,387),(374,388)),  
      11250 to 11280 => ((344,357),(345,359),(346,360),(373,387),(374,388),(375,389)),  
      11280 to 11310 => ((344,358),(345,359),(347,361),(374,388),(375,389),(376,390)),  
      11310 to 11340 => ((345,359),(346,360),(348,362),(375,389),(376,390),(377,391)),  
      11340 to 11370 => ((346,360),(347,361),(349,363),(376,390),(377,391),(378,392)),  
      11370 to 11400 => ((347,361),(348,362),(350,364),(377,391),(378,392),(379,393)),  
      11400 to 11430 => ((348,362),(349,363),(351,365),(378,392),(379,393),(380,394)),  
      11430 to 11460 => ((349,363),(350,364),(352,366),(379,393),(380,394),(381,395)),  
      11460 to 11490 => ((350,364),(351,365),(352,366),(380,394),(381,395),(382,396)),  
      11490 to 11520 => ((351,365),(352,366),(353,367),(381,395),(382,396),(383,397)),  
      11520 to 11550 => ((352,366),(353,367),(354,368),(382,396),(383,397),(384,398)),  
      11550 to 11580 => ((353,367),(354,368),(355,369),(383,397),(384,398),(386,400)),  
      11580 to 11610 => ((354,368),(355,369),(356,370),(384,398),(385,399),(387,401)),  
      11610 to 11640 => ((355,369),(356,370),(357,371),(385,399),(386,400),(388,402)),  
      11640 to 11670 => ((356,370),(357,371),(358,372),(386,400),(387,401),(389,403)),  
      11670 to 11700 => ((357,371),(358,372),(359,373),(387,401),(388,402),(390,404)),  
      11700 to 11730 => ((358,372),(359,373),(360,374),(388,402),(389,403),(391,405)),  
      11730 to 11760 => ((359,373),(360,374),(361,375),(389,403),(391,405),(392,406)),  
      11760 to 11790 => ((360,374),(361,375),(362,376),(390,404),(392,406),(393,407)),  
      11790 to 11820 => ((361,375),(362,376),(363,377),(391,405),(393,407),(394,408)),  
      11820 to 11850 => ((362,376),(363,377),(364,378),(392,406),(394,408),(395,409)),  
      11850 to 11880 => ((362,376),(364,378),(365,379),(393,407),(395,409),(396,410)),  
      11880 to 11910 => ((363,377),(365,379),(366,380),(394,408),(396,410),(397,411)),  
      11910 to 11940 => ((364,378),(366,380),(367,381),(395,409),(397,411),(398,412)),  
      11940 to 11970 => ((365,379),(367,381),(368,382),(396,410),(398,412),(399,413)),  
      11970 to 12000 => ((366,380),(368,382),(369,383),(398,412),(399,413),(400,414)),  
      12000 to 12030 => ((367,381),(369,383),(370,384),(399,413),(400,414),(401,415)),  
      12030 to 12060 => ((368,382),(370,384),(371,385),(400,414),(401,415),(402,416)),  
      12060 to 12090 => ((369,383),(370,384),(372,386),(401,415),(402,416),(403,417)),  
      12090 to 12120 => ((370,384),(371,385),(373,387),(402,416),(403,417),(404,418)),  
      12120 to 12150 => ((371,385),(372,386),(374,388),(403,417),(404,418),(405,419)),  
      12150 to 12180 => ((372,386),(373,387),(375,389),(404,418),(405,419),(406,420)),  
      12180 to 12210 => ((373,387),(374,388),(376,390),(405,419),(406,420),(407,421)),  
      12210 to 12250 => ((374,388),(375,389),(377,391),(406,420),(407,421),(408,422)),  
  );

 end package RoI_LUT_BOLA3;
