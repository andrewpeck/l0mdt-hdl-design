--------------------------------------------------------------------------------
--  UMass , Physics Department
--  Guillermo Loustau de Linares
--  gloustau@cern.ch
--------------------------------------------------------------------------------  
--  Project: ATLAS L0MDT Trigger 
--  Module: Hit Processor drift time and T0 compensation
--  Description:
--
--------------------------------------------------------------------------------
--  Revisions:
--      14/02/2019  0.1     File created
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;
use shared_lib.config_pkg.all;

package hps_rom_b_t0_pkg is
  -- integer values for T0 with 0.78 ns resolution
  -- T0 = ToF + t0
  -- t0 = 817 ; 542.5
  /*
  {"BIL", {{3, { 16.750000, 17.625000, 19.000000, 21.250000, 23.500000, 25.875000}}},},
  {"BML", {{3, { 24.125000, 25.500000, 27.875000, 30.875000, 33.500000, 36.750000}}},},
  {"BOL", {{3, { 32.000000, 33.750000, 36.500000, 40.125000, 44.875000, 49.500000}}},},
  */

  type t0LUT_chamber_t is array (0 to 7) of integer;
  type t0LUT_station_t is array (1 to 16) of t0LUT_chamber_t;
  
  constant c_BI_T0 : t0LUT_station_t :=(
    1  => (0,0,0,0,0,0,0,0), 
    2  => (0,0,0,0,0,0,0,0),
    3  => (716 , 717 , 719 , 722 , 724 , 728 , 0 , 0),
    4  => (0,0,0,0,0,0,0,0),
    5  => (0,0,0,0,0,0,0,0),
    6  => (0,0,0,0,0,0,0,0),
    7  => (0,0,0,0,0,0,0,0),
    8  => (0,0,0,0,0,0,0,0),
    9  => (0,0,0,0,0,0,0,0),
    10 => (0,0,0,0,0,0,0,0),
    11 => (0,0,0,0,0,0,0,0),
    12 => (0,0,0,0,0,0,0,0),
    13 => (0,0,0,0,0,0,0,0),
    14 => (0,0,0,0,0,0,0,0),
    15 => (0,0,0,0,0,0,0,0),
    16 => (0,0,0,0,0,0,0,0)
  );

  constant c_BM_T0 : t0LUT_station_t :=(
    1  => (0,0,0,0,0,0,0,0), 
    2  => (0,0,0,0,0,0,0,0),
    3  => (725 , 727 , 730 , 734 , 737 , 741 , 0 , 0 ),
    4  => (0,0,0,0,0,0,0,0),
    5  => (0,0,0,0,0,0,0,0),
    6  => (0,0,0,0,0,0,0,0),
    7  => (0,0,0,0,0,0,0,0),
    8  => (0,0,0,0,0,0,0,0),
    9  => (0,0,0,0,0,0,0,0),
    10 => (0,0,0,0,0,0,0,0),
    11 => (0,0,0,0,0,0,0,0),
    12 => (0,0,0,0,0,0,0,0),
    13 => (0,0,0,0,0,0,0,0),
    14 => (0,0,0,0,0,0,0,0),
    15 => (0,0,0,0,0,0,0,0),
    16 => (0,0,0,0,0,0,0,0)
  );

  constant c_BO_T0 : t0LUT_station_t :=(
    1  => (0,0,0,0,0,0,0,0), 
    2  => (0,0,0,0,0,0,0,0),
    3  => (735 , 738 , 741 , 746 , 752 , 758 , 0 , 0),
    4  => (0,0,0,0,0,0,0,0),
    5  => (0,0,0,0,0,0,0,0),
    6  => (0,0,0,0,0,0,0,0),
    7  => (0,0,0,0,0,0,0,0),
    8  => (0,0,0,0,0,0,0,0),
    9  => (0,0,0,0,0,0,0,0),
    10 => (0,0,0,0,0,0,0,0),
    11 => (0,0,0,0,0,0,0,0),
    12 => (0,0,0,0,0,0,0,0),
    13 => (0,0,0,0,0,0,0,0),
    14 => (0,0,0,0,0,0,0,0),
    15 => (0,0,0,0,0,0,0,0),
    16 => (0,0,0,0,0,0,0,0)
  );
    


    
end package hps_rom_b_t0_pkg;