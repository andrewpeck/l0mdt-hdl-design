--------------------------------------------------------------------------------
--  UMass , Physics Department
--  Guillermo Loustau de Linares
--  guillermo.ldl@cern.ch
--------------------------------------------------------------------------------  
--  Project: ATLAS L0MDT Trigger 
--  Module: PHI CENTER CHAMBER
--  Description: 
--
--------------------------------------------------------------------------------
--  Revisions:
--      2020.12.21  0.1     File created
--------------------------------------------------------------------------------


package mem_phi_center_chamber_pkg is
  
  
  
end package mem_phi_center_chamber_pkg;