library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;

package tar_pkg is

  constant TAR_PL_A_LATENCY : integer := 250;

end package tar_pkg;

------------------------------------------------------------

package body tar_pkg is

end package body tar_pkg;
