// SpyProtocol verilog include file.

// I chose these pretty arbitrarily. We can adjust as needed or add more
// valid metadata words.
parameter START_EVENT = 8'b10101011;
parameter END_EVENT = 8'b11001101;
