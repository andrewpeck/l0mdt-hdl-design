--------------------------------------------------------------------------------
--  UMass , Physics Department               
--  Yuan-Tang Chou                           
--  yuan-tang.chou@cern.ch                         
--------------------------------------------------------------------------------
--  Project: ATLAS L0MDT Trigger             
--  Module: Tube position coordinate 
--  Multiplier: 32 
--  Resolution: 0.03125 mm 
--  Description: Autogenerated file          
--                                           
--------------------------------------------------------------------------------
--  Revisions: 
--      
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package TC_B3A_pkg.vhd is
  constant MAX_TUBES_INN : 198;
  constant MAX_TUBES_MID : 296;
  constant MAX_TUBES_OUT : 400;
  -- constant MAX_TUBES_EXT : 5;
  type tube_coordinates_at is array (0 to 1) of real;
  type tube_coord_colum_aat is array (integer range <>) of tube_coordinates_at;
  type tube_coord_side_aat is array ( integer range <>) of tube_coord_colum_aat;    

  constant tube_coordinates_inn :  tube_coord_side_aat (0 to MAX_TUBES_INN - 1)(0 to 7):= (
    --     layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       , layer 6       , layer 7       ,
     0 => ((  330.017, 4770.928),(  315.000, 4796.938),(  330.017, 4822.950),(  315.000, 4848.961),(  315.000, 5048.998),(  330.017, 5075.009),(  315.000, 5101.020),(  330.017, 5127.031)), -- tube   0
     1 => ((  360.017, 4770.928),(  345.000, 4796.938),(  360.017, 4822.950),(  345.000, 4848.961),(  345.000, 5048.998),(  360.017, 5075.009),(  345.000, 5101.020),(  360.017, 5127.031)), -- tube   1
     2 => ((  390.052, 4770.928),(  375.035, 4796.938),(  390.052, 4822.950),(  375.035, 4848.961),(  375.035, 5048.998),(  390.052, 5075.009),(  375.035, 5101.020),(  390.052, 5127.031)), -- tube   2
     3 => ((  420.087, 4770.928),(  405.070, 4796.938),(  420.087, 4822.950),(  405.070, 4848.961),(  405.070, 5048.998),(  420.087, 5075.009),(  405.070, 5101.020),(  420.087, 5127.031)), -- tube   3
     4 => ((  450.122, 4770.928),(  435.105, 4796.938),(  450.122, 4822.950),(  435.105, 4848.961),(  435.105, 5048.998),(  450.122, 5075.009),(  435.105, 5101.020),(  450.122, 5127.031)), -- tube   4
     5 => ((  480.158, 4770.928),(  465.140, 4796.938),(  480.158, 4822.950),(  465.140, 4848.961),(  465.140, 5048.998),(  480.158, 5075.009),(  465.140, 5101.020),(  480.158, 5127.031)), -- tube   5
     6 => ((  510.193, 4770.928),(  495.175, 4796.938),(  510.193, 4822.950),(  495.175, 4848.961),(  495.175, 5048.998),(  510.193, 5075.009),(  495.175, 5101.020),(  510.193, 5127.031)), -- tube   6
     7 => ((  540.227, 4770.928),(  525.210, 4796.938),(  540.227, 4822.950),(  525.210, 4848.961),(  525.210, 5048.998),(  540.227, 5075.009),(  525.210, 5101.020),(  540.227, 5127.031)), -- tube   7
     8 => ((  570.263, 4770.928),(  555.245, 4796.938),(  570.263, 4822.950),(  555.245, 4848.961),(  555.245, 5048.998),(  570.263, 5075.009),(  555.245, 5101.020),(  570.263, 5127.031)), -- tube   8
     9 => ((  600.297, 4770.928),(  585.280, 4796.938),(  600.297, 4822.950),(  585.280, 4848.961),(  585.280, 5048.998),(  600.297, 5075.009),(  585.280, 5101.020),(  600.297, 5127.031)), -- tube   9
    10 => ((  630.333, 4770.928),(  615.315, 4796.938),(  630.333, 4822.950),(  615.315, 4848.961),(  615.315, 5048.998),(  630.333, 5075.009),(  615.315, 5101.020),(  630.333, 5127.031)), -- tube  10
    11 => ((  660.367, 4770.928),(  645.350, 4796.938),(  660.367, 4822.950),(  645.350, 4848.961),(  645.350, 5048.998),(  660.367, 5075.009),(  645.350, 5101.020),(  660.367, 5127.031)), -- tube  11
    12 => ((  690.403, 4770.928),(  675.385, 4796.938),(  690.438, 4822.950),(  675.420, 4848.961),(  675.385, 5048.998),(  690.403, 5075.009),(  675.385, 5101.020),(  690.403, 5127.031)), -- tube  12
    13 => ((  720.472, 4770.928),(  705.455, 4796.938),(  720.438, 4822.950),(  705.420, 4848.961),(  705.420, 5048.998),(  720.438, 5075.009),(  705.420, 5101.020),(  720.403, 5127.031)), -- tube  13
    14 => ((  750.472, 4770.928),(  735.455, 4796.938),(  750.472, 4822.950),(  735.455, 4848.961),(  735.455, 5048.998),(  750.472, 5075.009),(  735.455, 5101.020),(  750.508, 5127.031)), -- tube  14
    15 => ((  780.508, 4770.928),(  765.490, 4796.938),(  780.508, 4822.950),(  765.490, 4848.961),(  765.490, 5048.998),(  780.508, 5075.009),(  765.490, 5101.020),(  780.508, 5127.031)), -- tube  15
    16 => ((  810.542, 4770.928),(  795.525, 4796.938),(  810.542, 4822.950),(  795.525, 4848.961),(  795.525, 5048.998),(  810.542, 5075.009),(  795.525, 5101.020),(  810.508, 5127.031)), -- tube  16
    17 => ((  840.578, 4770.928),(  825.560, 4796.938),(  840.578, 4822.950),(  825.560, 4848.961),(  825.560, 5048.998),(  840.578, 5075.009),(  825.560, 5101.020),(  840.612, 5127.031)), -- tube  17
    18 => ((  870.612, 4770.928),(  855.595, 4796.938),(  870.612, 4822.950),(  855.595, 4848.961),(  855.595, 5048.998),(  870.612, 5075.009),(  855.595, 5101.020),(  870.612, 5127.031)), -- tube  18
    19 => ((  900.648, 4770.928),(  885.630, 4796.938),(  900.648, 4822.950),(  885.630, 4848.961),(  885.630, 5048.998),(  900.648, 5075.009),(  885.630, 5101.020),(  900.648, 5127.031)), -- tube  19
    20 => ((  930.682, 4770.928),(  915.665, 4796.938),(  930.682, 4822.950),(  915.665, 4848.961),(  915.665, 5048.998),(  930.648, 5075.009),(  915.665, 5101.020),(  930.682, 5127.031)), -- tube  20
    21 => ((  960.717, 4770.928),(  945.700, 4796.938),(  960.717, 4822.950),(  945.700, 4848.961),(  945.735, 5048.998),(  960.753, 5075.009),(  945.700, 5101.020),(  960.753, 5127.031)), -- tube  21
    22 => ((  990.753, 4770.928),(  975.735, 4796.938),(  990.753, 4822.950),(  975.735, 4848.961),(  975.735, 5048.998),(  990.753, 5075.009),(  975.735, 5101.020),(  990.753, 5127.031)), -- tube  22
    23 => (( 1020.787, 4770.928),( 1005.770, 4796.938),( 1020.787, 4822.950),( 1005.770, 4848.961),( 1005.770, 5048.998),( 1020.787, 5075.009),( 1005.805, 5101.020),( 1020.787, 5127.031)), -- tube  23
    24 => (( 1050.823, 4770.928),( 1035.805, 4796.938),( 1050.823, 4822.950),( 1035.805, 4848.961),( 1035.805, 5048.998),( 1050.823, 5075.009),( 1035.805, 5101.020),( 1050.823, 5127.031)), -- tube  24
    25 => (( 1080.858, 4770.928),( 1065.840, 4796.938),( 1080.858, 4822.950),( 1065.840, 4848.961),( 1065.840, 5048.998),( 1080.858, 5075.009),( 1065.840, 5101.020),( 1080.858, 5127.031)), -- tube  25
    26 => (( 1110.892, 4770.928),( 1095.875, 4796.938),( 1110.892, 4822.950),( 1095.875, 4848.961),( 1095.875, 5048.998),( 1110.892, 5075.009),( 1095.875, 5101.020),( 1110.892, 5127.031)), -- tube  26
    27 => (( 1140.927, 4770.928),( 1125.910, 4796.938),( 1140.927, 4822.950),( 1125.910, 4848.961),( 1125.910, 5048.998),( 1140.927, 5075.009),( 1125.910, 5101.020),( 1140.927, 5127.031)), -- tube  27
    28 => (( 1170.963, 4770.928),( 1155.945, 4796.938),( 1170.963, 4822.950),( 1155.945, 4848.961),( 1155.945, 5048.998),( 1170.963, 5075.009),( 1155.945, 5101.020),( 1170.963, 5127.031)), -- tube  28
    29 => (( 1200.997, 4770.928),( 1185.980, 4796.938),( 1200.997, 4822.950),( 1185.980, 4848.961),( 1185.980, 5048.998),( 1200.997, 5075.009),( 1185.980, 5101.020),( 1200.997, 5127.031)), -- tube  29
    30 => (( 1231.032, 4770.928),( 1216.015, 4796.938),( 1231.032, 4822.950),( 1216.015, 4848.961),( 1216.015, 5048.998),( 1231.032, 5075.009),( 1216.015, 5101.020),( 1231.032, 5127.031)), -- tube  30
    31 => (( 1280.017, 4770.928),( 1265.000, 4796.938),( 1280.017, 4822.950),( 1265.000, 4848.961),( 1265.000, 5048.998),( 1280.017, 5075.009),( 1265.000, 5101.020),( 1280.017, 5127.031)), -- tube  31
    32 => (( 1310.052, 4770.928),( 1295.035, 4796.938),( 1310.052, 4822.950),( 1295.035, 4848.961),( 1295.035, 5048.998),( 1310.052, 5075.009),( 1295.035, 5101.020),( 1310.052, 5127.031)), -- tube  32
    33 => (( 1340.088, 4770.928),( 1325.070, 4796.938),( 1340.088, 4822.950),( 1325.070, 4848.961),( 1325.070, 5048.998),( 1340.088, 5075.009),( 1325.070, 5101.020),( 1340.088, 5127.031)), -- tube  33
    34 => (( 1370.123, 4770.928),( 1355.105, 4796.938),( 1370.123, 4822.950),( 1355.105, 4848.961),( 1355.105, 5048.998),( 1370.123, 5075.009),( 1355.105, 5101.020),( 1370.123, 5127.031)), -- tube  34
    35 => (( 1400.157, 4770.928),( 1385.140, 4796.938),( 1400.157, 4822.950),( 1385.140, 4848.961),( 1385.140, 5048.998),( 1400.157, 5075.009),( 1385.140, 5101.020),( 1400.157, 5127.031)), -- tube  35
    36 => (( 1430.193, 4770.928),( 1415.175, 4796.938),( 1430.193, 4822.950),( 1415.175, 4848.961),( 1415.175, 5048.998),( 1430.193, 5075.009),( 1415.175, 5101.020),( 1430.193, 5127.031)), -- tube  36
    37 => (( 1460.228, 4770.928),( 1445.210, 4796.938),( 1460.228, 4822.950),( 1445.210, 4848.961),( 1445.210, 5048.998),( 1460.228, 5075.009),( 1445.210, 5101.020),( 1460.228, 5127.031)), -- tube  37
    38 => (( 1490.262, 4770.928),( 1475.245, 4796.938),( 1490.262, 4822.950),( 1475.245, 4848.961),( 1475.245, 5048.998),( 1490.262, 5075.009),( 1475.245, 5101.020),( 1490.262, 5127.031)), -- tube  38
    39 => (( 1520.297, 4770.928),( 1505.280, 4796.938),( 1520.297, 4822.950),( 1505.280, 4848.961),( 1505.280, 5048.998),( 1520.297, 5075.009),( 1505.280, 5101.020),( 1520.297, 5127.031)), -- tube  39
    40 => (( 1550.333, 4770.928),( 1535.315, 4796.938),( 1550.333, 4822.950),( 1535.315, 4848.961),( 1535.315, 5048.998),( 1550.333, 5075.009),( 1535.315, 5101.020),( 1550.333, 5127.031)), -- tube  40
    41 => (( 1580.368, 4770.928),( 1565.350, 4796.938),( 1580.368, 4822.950),( 1565.350, 4848.961),( 1565.350, 5048.998),( 1580.402, 5075.009),( 1565.350, 5101.020),( 1580.368, 5127.031)), -- tube  41
    42 => (( 1610.402, 4770.928),( 1595.385, 4796.938),( 1610.402, 4822.950),( 1595.385, 4848.961),( 1595.385, 5048.998),( 1610.402, 5075.009),( 1595.420, 5101.020),( 1610.402, 5127.031)), -- tube  42
    43 => (( 1640.438, 4770.928),( 1625.420, 4796.938),( 1640.438, 4822.950),( 1625.420, 4848.961),( 1625.420, 5048.998),( 1640.438, 5075.009),( 1625.420, 5101.020),( 1640.438, 5127.031)), -- tube  43
    44 => (( 1670.473, 4770.928),( 1655.455, 4796.938),( 1670.473, 4822.950),( 1655.455, 4848.961),( 1655.455, 5048.998),( 1670.473, 5075.009),( 1655.455, 5101.020),( 1670.473, 5127.031)), -- tube  44
    45 => (( 1700.507, 4770.928),( 1685.490, 4796.938),( 1700.507, 4822.950),( 1685.490, 4848.961),( 1685.490, 5048.998),( 1700.507, 5075.009),( 1685.490, 5101.020),( 1700.507, 5127.031)), -- tube  45
    46 => (( 1730.542, 4770.928),( 1715.525, 4796.938),( 1730.542, 4822.950),( 1715.525, 4848.961),( 1715.525, 5048.998),( 1730.542, 5075.009),( 1715.525, 5101.020),( 1730.542, 5127.031)), -- tube  46
    47 => (( 1760.578, 4770.928),( 1745.560, 4796.938),( 1760.578, 4822.950),( 1745.560, 4848.961),( 1745.560, 5048.998),( 1760.578, 5075.009),( 1745.560, 5101.020),( 1760.578, 5127.031)), -- tube  47
    48 => (( 1790.613, 4770.928),( 1775.595, 4796.938),( 1790.613, 4822.950),( 1775.595, 4848.961),( 1775.595, 5048.998),( 1790.613, 5075.009),( 1775.595, 5101.020),( 1790.613, 5127.031)), -- tube  48
    49 => (( 1820.647, 4770.928),( 1805.630, 4796.938),( 1820.647, 4822.950),( 1805.630, 4848.961),( 1805.630, 5048.998),( 1820.647, 5075.009),( 1805.630, 5101.020),( 1820.647, 5127.031)), -- tube  49
    50 => (( 1850.682, 4770.928),( 1835.665, 4796.938),( 1850.682, 4822.950),( 1835.665, 4848.961),( 1835.665, 5048.998),( 1850.682, 5075.009),( 1835.665, 5101.020),( 1850.682, 5127.031)), -- tube  50
    51 => (( 1880.718, 4770.928),( 1865.700, 4796.938),( 1880.718, 4822.950),( 1865.700, 4848.961),( 1865.700, 5048.998),( 1880.718, 5075.009),( 1865.700, 5101.020),( 1880.718, 5127.031)), -- tube  51
    52 => (( 1910.752, 4770.928),( 1895.735, 4796.938),( 1910.752, 4822.950),( 1895.735, 4848.961),( 1895.735, 5048.998),( 1910.752, 5075.009),( 1895.735, 5101.020),( 1910.752, 5127.031)), -- tube  52
    53 => (( 1940.787, 4770.928),( 1925.770, 4796.938),( 1940.787, 4822.950),( 1925.770, 4848.961),( 1925.770, 5048.998),( 1940.823, 5075.009),( 1925.770, 5101.020),( 1940.787, 5127.031)), -- tube  53
    54 => (( 1970.823, 4770.928),( 1955.805, 4796.938),( 1970.823, 4822.950),( 1955.805, 4848.961),( 1955.805, 5048.998),( 1970.823, 5075.009),( 1955.805, 5101.020),( 1970.823, 5127.031)), -- tube  54
    55 => (( 2000.858, 4770.928),( 1985.840, 4796.938),( 2000.858, 4822.950),( 1985.840, 4848.961),( 1985.840, 5048.998),( 2000.858, 5075.009),( 1985.840, 5101.020),( 2000.858, 5127.031)), -- tube  55
    56 => (( 2030.892, 4770.928),( 2015.875, 4796.938),( 2030.892, 4822.950),( 2015.875, 4848.961),( 2015.875, 5048.998),( 2030.892, 5075.009),( 2015.875, 5101.020),( 2030.892, 5127.031)), -- tube  56
    57 => (( 2060.927, 4770.928),( 2045.910, 4796.938),( 2060.927, 4822.950),( 2045.910, 4848.961),( 2045.910, 5048.998),( 2060.927, 5075.009),( 2045.910, 5101.020),( 2060.927, 5127.031)), -- tube  57
    58 => (( 2090.962, 4770.928),( 2075.945, 4796.938),( 2090.962, 4822.950),( 2075.945, 4848.961),( 2075.945, 5048.998),( 2090.962, 5075.009),( 2075.945, 5101.020),( 2090.962, 5127.031)), -- tube  58
    59 => (( 2120.998, 4770.928),( 2105.980, 4796.938),( 2120.998, 4822.950),( 2105.980, 4848.961),( 2105.980, 5048.998),( 2120.998, 5075.009),( 2105.980, 5101.020),( 2120.998, 5127.031)), -- tube  59
    60 => (( 2151.067, 4770.928),( 2136.015, 4796.938),( 2151.032, 4822.950),( 2136.015, 4848.961),( 2136.015, 5048.998),( 2151.032, 5075.009),( 2136.015, 5101.020),( 2151.032, 5127.031)), -- tube  60
    61 => (( 2181.067, 4770.928),( 2166.050, 4796.938),( 2181.067, 4822.950),( 2166.050, 4848.961),( 2166.050, 5048.998),( 2181.067, 5075.009),( 2166.050, 5101.020),( 2181.067, 5127.031)), -- tube  61
    62 => (( 2211.103, 4770.928),( 2196.085, 4796.938),( 2211.103, 4822.950),( 2196.085, 4848.961),( 2196.085, 5048.998),( 2211.103, 5075.009),( 2196.085, 5101.020),( 2211.103, 5127.031)), -- tube  62
    63 => (( 2241.137, 4770.928),( 2226.120, 4796.938),( 2241.137, 4822.950),( 2226.120, 4848.961),( 2226.120, 5048.998),( 2241.137, 5075.009),( 2226.120, 5101.020),( 2241.137, 5127.031)), -- tube  63
    64 => (( 2271.173, 4770.928),( 2256.155, 4796.938),( 2271.173, 4822.950),( 2256.155, 4848.961),( 2256.155, 5048.998),( 2271.173, 5075.009),( 2256.155, 5101.020),( 2271.173, 5127.031)), -- tube  64
    65 => (( 2301.242, 4770.928),( 2286.190, 4796.938),( 2301.208, 4822.950),( 2286.190, 4848.961),( 2286.190, 5048.998),( 2301.208, 5075.009),( 2286.190, 5101.020),( 2301.208, 5127.031)), -- tube  65
    66 => (( 2331.242, 4770.928),( 2316.225, 4796.938),( 2331.242, 4822.950),( 2316.225, 4848.961),( 2316.225, 5048.998),( 2331.242, 5075.009),( 2316.225, 5101.020),( 2331.242, 5127.031)), -- tube  66
    67 => (( 2380.018, 4770.928),( 2365.000, 4796.938),( 2380.052, 4822.950),( 2365.000, 4848.961),( 2365.000, 5048.998),( 2380.018, 5075.009),( 2365.000, 5101.020),( 2380.018, 5127.031)), -- tube  67
    68 => (( 2410.052, 4770.928),( 2395.035, 4796.938),( 2410.052, 4822.950),( 2395.035, 4848.961),( 2395.035, 5048.998),( 2410.052, 5075.009),( 2395.035, 5101.020),( 2410.052, 5127.031)), -- tube  68
    69 => (( 2440.087, 4770.928),( 2425.070, 4796.938),( 2440.087, 4822.950),( 2425.070, 4848.961),( 2425.070, 5048.998),( 2440.087, 5075.009),( 2425.070, 5101.020),( 2440.087, 5127.031)), -- tube  69
    70 => (( 2470.123, 4770.928),( 2455.105, 4796.938),( 2470.123, 4822.950),( 2455.105, 4848.961),( 2455.105, 5048.998),( 2470.123, 5075.009),( 2455.105, 5101.020),( 2470.123, 5127.031)), -- tube  70
    71 => (( 2500.157, 4770.928),( 2485.140, 4796.938),( 2500.157, 4822.950),( 2485.140, 4848.961),( 2485.140, 5048.998),( 2500.157, 5075.009),( 2485.140, 5101.020),( 2500.157, 5127.031)), -- tube  71
    72 => (( 2530.192, 4770.928),( 2515.175, 4796.938),( 2530.192, 4822.950),( 2515.175, 4848.961),( 2515.175, 5048.998),( 2530.192, 5075.009),( 2515.175, 5101.020),( 2530.192, 5127.031)), -- tube  72
    73 => (( 2560.228, 4770.928),( 2545.210, 4796.938),( 2560.228, 4822.950),( 2545.210, 4848.961),( 2545.210, 5048.998),( 2560.228, 5075.009),( 2545.210, 5101.020),( 2560.228, 5127.031)), -- tube  73
    74 => (( 2590.262, 4770.928),( 2575.245, 4796.938),( 2590.262, 4822.950),( 2575.245, 4848.961),( 2575.245, 5048.998),( 2590.262, 5075.009),( 2575.245, 5101.020),( 2590.262, 5127.031)), -- tube  74
    75 => (( 2620.298, 4770.928),( 2605.280, 4796.938),( 2620.298, 4822.950),( 2605.280, 4848.961),( 2605.280, 5048.998),( 2620.298, 5075.009),( 2605.280, 5101.020),( 2620.298, 5127.031)), -- tube  75
    76 => (( 2650.333, 4770.928),( 2635.315, 4796.938),( 2650.333, 4822.950),( 2635.315, 4848.961),( 2635.315, 5048.998),( 2650.333, 5075.009),( 2635.315, 5101.020),( 2650.333, 5127.031)), -- tube  76
    77 => (( 2680.367, 4770.928),( 2665.350, 4796.938),( 2680.367, 4822.950),( 2665.350, 4848.961),( 2665.350, 5048.998),( 2680.367, 5075.009),( 2665.350, 5101.020),( 2680.367, 5127.031)), -- tube  77
    78 => (( 2710.403, 4770.928),( 2695.385, 4796.938),( 2710.403, 4822.950),( 2695.385, 4848.961),( 2695.385, 5048.998),( 2710.403, 5075.009),( 2695.385, 5101.020),( 2710.403, 5127.031)), -- tube  78
    79 => (( 2740.438, 4770.928),( 2725.420, 4796.938),( 2740.438, 4822.950),( 2725.420, 4848.961),( 2725.420, 5048.998),( 2740.438, 5075.009),( 2725.420, 5101.020),( 2740.438, 5127.031)), -- tube  79
    80 => (( 2770.472, 4770.928),( 2755.455, 4796.938),( 2770.472, 4822.950),( 2755.455, 4848.961),( 2755.455, 5048.998),( 2770.472, 5075.009),( 2755.455, 5101.020),( 2770.472, 5127.031)), -- tube  80
    81 => (( 2800.508, 4770.928),( 2785.490, 4796.938),( 2800.508, 4822.950),( 2785.490, 4848.961),( 2785.490, 5048.998),( 2800.508, 5075.009),( 2785.490, 5101.020),( 2800.508, 5127.031)), -- tube  81
    82 => (( 2830.542, 4770.928),( 2815.525, 4796.938),( 2830.542, 4822.950),( 2815.525, 4848.961),( 2815.525, 5048.998),( 2830.542, 5075.009),( 2815.525, 5101.020),( 2830.542, 5127.031)), -- tube  82
    83 => (( 2860.577, 4770.928),( 2845.560, 4796.938),( 2860.577, 4822.950),( 2845.560, 4848.961),( 2845.560, 5048.998),( 2860.577, 5075.009),( 2845.560, 5101.020),( 2860.577, 5127.031)), -- tube  83
    84 => (( 2890.613, 4770.928),( 2875.595, 4796.938),( 2890.613, 4822.950),( 2875.595, 4848.961),( 2875.595, 5048.998),( 2890.613, 5075.009),( 2875.595, 5101.020),( 2890.613, 5127.031)), -- tube  84
    85 => (( 2920.647, 4770.928),( 2905.630, 4796.938),( 2920.647, 4822.950),( 2905.630, 4848.961),( 2905.630, 5048.998),( 2920.647, 5075.009),( 2905.630, 5101.020),( 2920.647, 5127.031)), -- tube  85
    86 => (( 2950.683, 4770.928),( 2935.665, 4796.938),( 2950.683, 4822.950),( 2935.665, 4848.961),( 2935.665, 5048.998),( 2950.683, 5075.009),( 2935.665, 5101.020),( 2950.683, 5127.031)), -- tube  86
    87 => (( 2980.718, 4770.928),( 2965.700, 4796.938),( 2980.718, 4822.950),( 2965.700, 4848.961),( 2965.700, 5048.998),( 2980.718, 5075.009),( 2965.700, 5101.020),( 2980.718, 5127.031)), -- tube  87
    88 => (( 3010.752, 4770.928),( 2995.735, 4796.938),( 3010.752, 4822.950),( 2995.735, 4848.961),( 2995.735, 5048.998),( 3010.752, 5075.009),( 2995.735, 5101.020),( 3010.752, 5127.031)), -- tube  88
    89 => (( 3040.788, 4770.928),( 3025.770, 4796.938),( 3040.788, 4822.950),( 3025.770, 4848.961),( 3025.770, 5048.998),( 3040.788, 5075.009),( 3025.770, 5101.020),( 3040.788, 5127.031)), -- tube  89
    90 => (( 3070.823, 4770.928),( 3055.805, 4796.938),( 3070.823, 4822.950),( 3055.805, 4848.961),( 3055.805, 5048.998),( 3070.823, 5075.009),( 3055.805, 5101.020),( 3070.823, 5127.031)), -- tube  90
    91 => (( 3100.857, 4770.928),( 3085.840, 4796.938),( 3100.857, 4822.950),( 3085.840, 4848.961),( 3085.840, 5048.998),( 3100.857, 5075.009),( 3085.840, 5101.020),( 3100.857, 5127.031)), -- tube  91
    92 => (( 3130.893, 4770.928),( 3115.875, 4796.938),( 3130.893, 4822.950),( 3115.875, 4848.961),( 3115.875, 5048.998),( 3130.893, 5075.009),( 3115.875, 5101.020),( 3130.893, 5127.031)), -- tube  92
    93 => (( 3160.927, 4770.928),( 3145.910, 4796.938),( 3160.927, 4822.950),( 3145.910, 4848.961),( 3145.910, 5048.998),( 3160.927, 5075.009),( 3145.910, 5101.020),( 3160.927, 5127.031)), -- tube  93
    94 => (( 3190.962, 4770.928),( 3175.945, 4796.938),( 3190.962, 4822.950),( 3175.945, 4848.961),( 3175.945, 5048.998),( 3190.962, 5075.009),( 3175.945, 5101.020),( 3190.962, 5127.031)), -- tube  94
    95 => (( 3220.998, 4770.928),( 3205.980, 4796.938),( 3220.998, 4822.950),( 3205.980, 4848.961),( 3205.980, 5048.998),( 3220.998, 5075.009),( 3205.980, 5101.020),( 3220.998, 5127.031)), -- tube  95
    96 => (( 3251.032, 4770.928),( 3236.015, 4796.938),( 3251.032, 4822.950),( 3236.015, 4848.961),( 3236.015, 5048.998),( 3251.032, 5075.009),( 3236.015, 5101.020),( 3251.032, 5127.031)), -- tube  96
    97 => (( 3480.018, 4770.928),( 3465.000, 4796.938),( 3480.018, 4822.950),( 3465.000, 4848.961),( 3465.000, 5048.998),( 3480.018, 5075.009),( 3465.035, 5101.020),( 3480.018, 5127.031)), -- tube  97
    98 => (( 3510.052, 4770.928),( 3495.035, 4796.938),( 3510.052, 4822.950),( 3495.035, 4848.961),( 3495.035, 5048.998),( 3510.052, 5075.009),( 3495.035, 5101.020),( 3510.052, 5127.031)), -- tube  98
    99 => (( 3540.087, 4770.928),( 3525.070, 4796.938),( 3540.087, 4822.950),( 3525.070, 4848.961),( 3525.070, 5048.998),( 3540.087, 5075.009),( 3525.070, 5101.020),( 3540.087, 5127.031)), -- tube  99
   100 => (( 3570.123, 4770.928),( 3555.105, 4796.938),( 3570.123, 4822.950),( 3555.105, 4848.961),( 3555.105, 5048.998),( 3570.123, 5075.009),( 3555.105, 5101.020),( 3570.123, 5127.031)), -- tube 100
   101 => (( 3600.157, 4770.928),( 3585.140, 4796.938),( 3600.157, 4822.950),( 3585.140, 4848.961),( 3585.140, 5048.998),( 3600.157, 5075.009),( 3585.140, 5101.020),( 3600.157, 5127.031)), -- tube 101
   102 => (( 3630.192, 4770.928),( 3615.175, 4796.938),( 3630.192, 4822.950),( 3615.175, 4848.961),( 3615.175, 5048.998),( 3630.228, 5075.009),( 3615.175, 5101.020),( 3630.192, 5127.031)), -- tube 102
   103 => (( 3660.228, 4770.928),( 3645.210, 4796.938),( 3660.228, 4822.950),( 3645.210, 4848.961),( 3645.210, 5048.998),( 3660.228, 5075.009),( 3645.210, 5101.020),( 3660.228, 5127.031)), -- tube 103
   104 => (( 3690.262, 4770.928),( 3675.245, 4796.938),( 3690.262, 4822.950),( 3675.245, 4848.961),( 3675.245, 5048.998),( 3690.262, 5075.009),( 3675.245, 5101.020),( 3690.262, 5127.031)), -- tube 104
   105 => (( 3720.298, 4770.928),( 3705.280, 4796.938),( 3720.298, 4822.950),( 3705.280, 4848.961),( 3705.280, 5048.998),( 3720.298, 5075.009),( 3705.280, 5101.020),( 3720.298, 5127.031)), -- tube 105
   106 => (( 3750.333, 4770.928),( 3735.315, 4796.938),( 3750.333, 4822.950),( 3735.315, 4848.961),( 3735.315, 5048.998),( 3750.333, 5075.009),( 3735.315, 5101.020),( 3750.333, 5127.031)), -- tube 106
   107 => (( 3780.367, 4770.928),( 3765.350, 4796.938),( 3780.367, 4822.950),( 3765.350, 4848.961),( 3765.350, 5048.998),( 3780.367, 5075.009),( 3765.350, 5101.020),( 3780.367, 5127.031)), -- tube 107
   108 => (( 3810.403, 4770.928),( 3795.385, 4796.938),( 3810.438, 4822.950),( 3795.385, 4848.961),( 3795.385, 5048.998),( 3810.403, 5075.009),( 3795.385, 5101.020),( 3810.403, 5127.031)), -- tube 108
   109 => (( 3840.438, 4770.928),( 3825.420, 4796.938),( 3840.438, 4822.950),( 3825.420, 4848.961),( 3825.420, 5048.998),( 3840.438, 5075.009),( 3825.420, 5101.020),( 3840.438, 5127.031)), -- tube 109
   110 => (( 3870.472, 4770.928),( 3855.455, 4796.938),( 3870.472, 4822.950),( 3855.455, 4848.961),( 3855.455, 5048.998),( 3870.472, 5075.009),( 3855.455, 5101.020),( 3870.472, 5127.031)), -- tube 110
   111 => (( 3900.508, 4770.928),( 3885.490, 4796.938),( 3900.508, 4822.950),( 3885.490, 4848.961),( 3885.490, 5048.998),( 3900.508, 5075.009),( 3885.490, 5101.020),( 3900.508, 5127.031)), -- tube 111
   112 => (( 3930.542, 4770.928),( 3915.525, 4796.938),( 3930.542, 4822.950),( 3915.525, 4848.961),( 3915.525, 5048.998),( 3930.542, 5075.009),( 3915.525, 5101.020),( 3930.542, 5127.031)), -- tube 112
   113 => (( 3960.577, 4770.928),( 3945.560, 4796.938),( 3960.577, 4822.950),( 3945.560, 4848.961),( 3945.560, 5048.998),( 3960.577, 5075.009),( 3945.560, 5101.020),( 3960.577, 5127.031)), -- tube 113
   114 => (( 3990.613, 4770.928),( 3975.595, 4796.938),( 3990.613, 4822.950),( 3975.595, 4848.961),( 3975.595, 5048.998),( 3990.613, 5075.009),( 3975.595, 5101.020),( 3990.613, 5127.031)), -- tube 114
   115 => (( 4020.647, 4770.928),( 4005.630, 4796.938),( 4020.647, 4822.950),( 4005.630, 4848.961),( 4005.630, 5048.998),( 4020.647, 5075.009),( 4005.630, 5101.020),( 4020.647, 5127.031)), -- tube 115
   116 => (( 4050.683, 4770.928),( 4035.665, 4796.938),( 4050.683, 4822.950),( 4035.665, 4848.961),( 4035.665, 5048.998),( 4050.683, 5075.009),( 4035.665, 5101.020),( 4050.683, 5127.031)), -- tube 116
   117 => (( 4080.718, 4770.928),( 4065.700, 4796.938),( 4080.718, 4822.950),( 4065.700, 4848.961),( 4065.700, 5048.998),( 4080.718, 5075.009),( 4065.700, 5101.020),( 4080.718, 5127.031)), -- tube 117
   118 => (( 4110.752, 4770.928),( 4095.735, 4796.938),( 4110.752, 4822.950),( 4095.735, 4848.961),( 4095.735, 5048.998),( 4110.752, 5075.009),( 4095.735, 5101.020),( 4110.752, 5127.031)), -- tube 118
   119 => (( 4140.788, 4770.928),( 4125.770, 4796.938),( 4140.788, 4822.950),( 4125.770, 4848.961),( 4125.770, 5048.998),( 4140.788, 5075.009),( 4125.770, 5101.020),( 4140.788, 5127.031)), -- tube 119
   120 => (( 4170.822, 4770.928),( 4155.805, 4796.938),( 4170.822, 4822.950),( 4155.805, 4848.961),( 4155.805, 5048.998),( 4170.822, 5075.009),( 4155.805, 5101.020),( 4170.822, 5127.031)), -- tube 120
   121 => (( 4200.857, 4770.928),( 4185.840, 4796.938),( 4200.857, 4822.950),( 4185.840, 4848.961),( 4185.840, 5048.998),( 4200.857, 5075.009),( 4185.840, 5101.020),( 4200.857, 5127.031)), -- tube 121
   122 => (( 4230.893, 4770.928),( 4215.875, 4796.938),( 4230.893, 4822.950),( 4215.875, 4848.961),( 4215.875, 5048.998),( 4230.893, 5075.009),( 4215.875, 5101.020),( 4230.893, 5127.031)), -- tube 122
   123 => (( 4260.928, 4770.928),( 4245.910, 4796.938),( 4260.928, 4822.950),( 4245.910, 4848.961),( 4245.910, 5048.998),( 4260.928, 5075.009),( 4245.910, 5101.020),( 4260.928, 5127.031)), -- tube 123
   124 => (( 4290.962, 4770.928),( 4275.945, 4796.938),( 4290.962, 4822.950),( 4275.945, 4848.961),( 4275.945, 5048.998),( 4290.962, 5075.009),( 4275.945, 5101.020),( 4290.962, 5127.031)), -- tube 124
   125 => (( 4320.998, 4770.928),( 4305.980, 4796.938),( 4320.998, 4822.950),( 4305.980, 4848.961),( 4305.980, 5048.998),( 4320.998, 5075.009),( 4305.980, 5101.020),( 4320.998, 5127.031)), -- tube 125
   126 => (( 4351.033, 4770.928),( 4336.015, 4796.938),( 4351.033, 4822.950),( 4336.015, 4848.961),( 4336.015, 5048.998),( 4351.033, 5075.009),( 4336.015, 5101.020),( 4351.033, 5127.031)), -- tube 126
   127 => (( 4381.067, 4770.928),( 4366.050, 4796.938),( 4381.067, 4822.950),( 4366.050, 4848.961),( 4366.050, 5048.998),( 4381.067, 5075.009),( 4366.050, 5101.020),( 4381.067, 5127.031)), -- tube 127
   128 => (( 4411.103, 4770.928),( 4396.085, 4796.938),( 4411.103, 4822.950),( 4396.085, 4848.961),( 4396.085, 5048.998),( 4411.103, 5075.009),( 4396.085, 5101.020),( 4411.103, 5127.031)), -- tube 128
   129 => (( 4441.138, 4770.928),( 4426.120, 4796.938),( 4441.138, 4822.950),( 4426.120, 4848.961),( 4426.120, 5048.998),( 4441.138, 5075.009),( 4426.120, 5101.020),( 4441.138, 5127.031)), -- tube 129
   130 => (( 4471.172, 4770.928),( 4456.155, 4796.938),( 4471.172, 4822.950),( 4456.155, 4848.961),( 4456.155, 5048.998),( 4471.172, 5075.009),( 4456.155, 5101.020),( 4471.172, 5127.031)), -- tube 130
   131 => (( 4501.208, 4770.928),( 4486.190, 4796.938),( 4501.208, 4822.950),( 4486.190, 4848.961),( 4486.190, 5048.998),( 4501.208, 5075.009),( 4486.190, 5101.020),( 4501.208, 5127.031)), -- tube 131
   132 => (( 4531.243, 4770.928),( 4516.225, 4796.938),( 4531.243, 4822.950),( 4516.225, 4848.961),( 4516.225, 5048.998),( 4531.243, 5075.009),( 4516.225, 5101.020),( 4531.243, 5127.031)), -- tube 132
   133 => (( 4580.018, 4770.928),( 4565.000, 4796.938),( 4580.018, 4822.950),( 4565.000, 4848.961),( 4565.000, 5048.998),( 4580.018, 5075.009),( 4565.000, 5101.020),( 4580.018, 5127.031)), -- tube 133
   134 => (( 4610.053, 4770.928),( 4595.035, 4796.938),( 4610.053, 4822.950),( 4595.035, 4848.961),( 4595.035, 5048.998),( 4610.053, 5075.009),( 4595.035, 5101.020),( 4610.053, 5127.031)), -- tube 134
   135 => (( 4640.087, 4770.928),( 4625.070, 4796.938),( 4640.087, 4822.950),( 4625.070, 4848.961),( 4625.070, 5048.998),( 4640.087, 5075.009),( 4625.070, 5101.020),( 4640.087, 5127.031)), -- tube 135
   136 => (( 4670.123, 4770.928),( 4655.105, 4796.938),( 4670.123, 4822.950),( 4655.105, 4848.961),( 4655.105, 5048.998),( 4670.123, 5075.009),( 4655.105, 5101.020),( 4670.123, 5127.031)), -- tube 136
   137 => (( 4700.158, 4770.928),( 4685.140, 4796.938),( 4700.158, 4822.950),( 4685.140, 4848.961),( 4685.140, 5048.998),( 4700.158, 5075.009),( 4685.140, 5101.020),( 4700.158, 5127.031)), -- tube 137
   138 => (( 4730.192, 4770.928),( 4715.175, 4796.938),( 4730.192, 4822.950),( 4715.175, 4848.961),( 4715.175, 5048.998),( 4730.192, 5075.009),( 4715.175, 5101.020),( 4730.192, 5127.031)), -- tube 138
   139 => (( 4760.228, 4770.928),( 4745.210, 4796.938),( 4760.228, 4822.950),( 4745.210, 4848.961),( 4745.210, 5048.998),( 4760.228, 5075.009),( 4745.210, 5101.020),( 4760.228, 5127.031)), -- tube 139
   140 => (( 4790.263, 4770.928),( 4775.245, 4796.938),( 4790.263, 4822.950),( 4775.245, 4848.961),( 4775.245, 5048.998),( 4790.263, 5075.009),( 4775.245, 5101.020),( 4790.263, 5127.031)), -- tube 140
   141 => (( 4820.297, 4770.928),( 4805.280, 4796.938),( 4820.297, 4822.950),( 4805.280, 4848.961),( 4805.280, 5048.998),( 4820.297, 5075.009),( 4805.280, 5101.020),( 4820.297, 5127.031)), -- tube 141
   142 => (( 4850.333, 4770.928),( 4835.315, 4796.938),( 4850.333, 4822.950),( 4835.315, 4848.961),( 4835.315, 5048.998),( 4850.333, 5075.009),( 4835.315, 5101.020),( 4850.333, 5127.031)), -- tube 142
   143 => (( 4880.368, 4770.928),( 4865.350, 4796.938),( 4880.368, 4822.950),( 4865.350, 4848.961),( 4865.350, 5048.998),( 4880.368, 5075.009),( 4865.350, 5101.020),( 4880.368, 5127.031)), -- tube 143
   144 => (( 4910.402, 4770.928),( 4895.385, 4796.938),( 4910.402, 4822.950),( 4895.385, 4848.961),( 4895.385, 5048.998),( 4910.402, 5075.009),( 4895.385, 5101.020),( 4910.402, 5127.031)), -- tube 144
   145 => (( 4940.438, 4770.928),( 4925.420, 4796.938),( 4940.438, 4822.950),( 4925.420, 4848.961),( 4925.420, 5048.998),( 4940.438, 5075.009),( 4925.420, 5101.020),( 4940.438, 5127.031)), -- tube 145
   146 => (( 4970.473, 4770.928),( 4955.455, 4796.938),( 4970.473, 4822.950),( 4955.455, 4848.961),( 4955.455, 5048.998),( 4970.473, 5075.009),( 4955.455, 5101.020),( 4970.473, 5127.031)), -- tube 146
   147 => (( 5000.507, 4770.928),( 4985.490, 4796.938),( 5000.507, 4822.950),( 4985.490, 4848.961),( 4985.490, 5048.998),( 5000.507, 5075.009),( 4985.490, 5101.020),( 5000.507, 5127.031)), -- tube 147
   148 => (( 5030.542, 4770.928),( 5015.525, 4796.938),( 5030.542, 4822.950),( 5015.525, 4848.961),( 5015.525, 5048.998),( 5030.542, 5075.009),( 5015.525, 5101.020),( 5030.542, 5127.031)), -- tube 148
   149 => (( 5060.578, 4770.928),( 5045.560, 4796.938),( 5060.578, 4822.950),( 5045.560, 4848.961),( 5045.560, 5048.998),( 5060.578, 5075.009),( 5045.560, 5101.020),( 5060.578, 5127.031)), -- tube 149
   150 => (( 5090.612, 4770.928),( 5075.595, 4796.938),( 5090.612, 4822.950),( 5075.595, 4848.961),( 5075.595, 5048.998),( 5090.612, 5075.009),( 5075.595, 5101.020),( 5090.612, 5127.031)), -- tube 150
   151 => (( 5120.647, 4770.928),( 5105.630, 4796.938),( 5120.647, 4822.950),( 5105.630, 4848.961),( 5105.630, 5048.998),( 5120.647, 5075.009),( 5105.630, 5101.020),( 5120.647, 5127.031)), -- tube 151
   152 => (( 5150.683, 4770.928),( 5135.665, 4796.938),( 5150.683, 4822.950),( 5135.665, 4848.961),( 5135.665, 5048.998),( 5150.683, 5075.009),( 5135.665, 5101.020),( 5150.683, 5127.031)), -- tube 152
   153 => (( 5180.717, 4770.928),( 5165.700, 4796.938),( 5180.717, 4822.950),( 5165.700, 4848.961),( 5165.700, 5048.998),( 5180.717, 5075.009),( 5165.700, 5101.020),( 5180.717, 5127.031)), -- tube 153
   154 => (( 5210.752, 4770.928),( 5195.735, 4796.938),( 5210.752, 4822.950),( 5195.735, 4848.961),( 5195.735, 5048.998),( 5210.752, 5075.009),( 5195.735, 5101.020),( 5210.752, 5127.031)), -- tube 154
   155 => (( 5240.788, 4770.928),( 5225.770, 4796.938),( 5240.788, 4822.950),( 5225.770, 4848.961),( 5225.770, 5048.998),( 5240.788, 5075.009),( 5225.770, 5101.020),( 5240.788, 5127.031)), -- tube 155
   156 => (( 5270.822, 4770.928),( 5255.805, 4796.938),( 5270.822, 4822.950),( 5255.805, 4848.961),( 5255.805, 5048.998),( 5270.822, 5075.009),( 5255.805, 5101.020),( 5270.822, 5127.031)), -- tube 156
   157 => (( 5300.857, 4770.928),( 5285.840, 4796.938),( 5300.857, 4822.950),( 5285.840, 4848.961),( 5285.840, 5048.998),( 5300.857, 5075.009),( 5285.840, 5101.020),( 5300.857, 5127.031)), -- tube 157
   158 => (( 5330.893, 4770.928),( 5315.875, 4796.938),( 5330.893, 4822.950),( 5315.875, 4848.961),( 5315.875, 5048.998),( 5330.893, 5075.009),( 5315.875, 5101.020),( 5330.893, 5127.031)), -- tube 158
   159 => (( 5360.928, 4770.928),( 5345.910, 4796.938),( 5360.928, 4822.950),( 5345.910, 4848.961),( 5345.910, 5048.998),( 5360.928, 5075.009),( 5345.910, 5101.020),( 5360.928, 5127.031)), -- tube 159
   160 => (( 5390.962, 4770.928),( 5375.945, 4796.938),( 5390.962, 4822.950),( 5375.945, 4848.961),( 5375.945, 5048.998),( 5390.962, 5075.009),( 5375.945, 5101.020),( 5390.962, 5127.031)), -- tube 160
   161 => (( 5420.998, 4770.928),( 5405.980, 4796.938),( 5420.998, 4822.950),( 5405.980, 4848.961),( 5405.980, 5048.998),( 5420.998, 5075.009),( 5405.980, 5101.020),( 5420.998, 5127.031)), -- tube 161
   162 => (( 5451.033, 4770.928),( 5436.015, 4796.938),( 5451.033, 4822.950),( 5436.015, 4848.961),( 5436.015, 5048.998),( 5451.033, 5075.009),( 5436.015, 5101.020),( 5451.033, 5127.031)), -- tube 162
   163 => (( 5500.018, 4770.928),( 5485.000, 4796.938),( 5500.018, 4822.950),( 5485.000, 4848.961),( 5485.000, 5048.998),( 5500.018, 5075.009),( 5485.000, 5101.020),( 5500.018, 5127.031)), -- tube 163
   164 => (( 5530.053, 4770.928),( 5515.035, 4796.938),( 5530.053, 4822.950),( 5515.035, 4848.961),( 5515.035, 5048.998),( 5530.053, 5075.009),( 5515.035, 5101.020),( 5530.053, 5127.031)), -- tube 164
   165 => (( 5560.087, 4770.928),( 5545.070, 4796.938),( 5560.087, 4822.950),( 5545.070, 4848.961),( 5545.070, 5048.998),( 5560.087, 5075.009),( 5545.070, 5101.020),( 5560.087, 5127.031)), -- tube 165
   166 => (( 5590.123, 4770.928),( 5575.105, 4796.938),( 5590.123, 4822.950),( 5575.105, 4848.961),( 5575.105, 5048.998),( 5590.123, 5075.009),( 5575.105, 5101.020),( 5590.123, 5127.031)), -- tube 166
   167 => (( 5620.158, 4770.928),( 5605.140, 4796.938),( 5620.158, 4822.950),( 5605.140, 4848.961),( 5605.140, 5048.998),( 5620.158, 5075.009),( 5605.140, 5101.020),( 5620.158, 5127.031)), -- tube 167
   168 => (( 5650.192, 4770.928),( 5635.175, 4796.938),( 5650.192, 4822.950),( 5635.175, 4848.961),( 5635.175, 5048.998),( 5650.192, 5075.009),( 5635.175, 5101.020),( 5650.192, 5127.031)), -- tube 168
   169 => (( 5680.228, 4770.928),( 5665.210, 4796.938),( 5680.228, 4822.950),( 5665.210, 4848.961),( 5665.210, 5048.998),( 5680.228, 5075.009),( 5665.210, 5101.020),( 5680.228, 5127.031)), -- tube 169
   170 => (( 5710.263, 4770.928),( 5695.245, 4796.938),( 5710.263, 4822.950),( 5695.245, 4848.961),( 5695.245, 5048.998),( 5710.263, 5075.009),( 5695.245, 5101.020),( 5710.263, 5127.031)), -- tube 170
   171 => (( 5740.297, 4770.928),( 5725.280, 4796.938),( 5740.297, 4822.950),( 5725.280, 4848.961),( 5725.280, 5048.998),( 5740.297, 5075.009),( 5725.280, 5101.020),( 5740.297, 5127.031)), -- tube 171
   172 => (( 5770.333, 4770.928),( 5755.315, 4796.938),( 5770.333, 4822.950),( 5755.315, 4848.961),( 5755.315, 5048.998),( 5770.333, 5075.009),( 5755.315, 5101.020),( 5770.333, 5127.031)), -- tube 172
   173 => (( 5800.368, 4770.928),( 5785.350, 4796.938),( 5800.368, 4822.950),( 5785.350, 4848.961),( 5785.350, 5048.998),( 5800.368, 5075.009),( 5785.350, 5101.020),( 5800.368, 5127.031)), -- tube 173
   174 => (( 5830.402, 4770.928),( 5815.385, 4796.938),( 5830.402, 4822.950),( 5815.385, 4848.961),( 5815.385, 5048.998),( 5830.402, 5075.009),( 5815.385, 5101.020),( 5830.402, 5127.031)), -- tube 174
   175 => (( 5860.438, 4770.928),( 5845.420, 4796.938),( 5860.438, 4822.950),( 5845.420, 4848.961),( 5845.420, 5048.998),( 5860.438, 5075.009),( 5845.420, 5101.020),( 5860.438, 5127.031)), -- tube 175
   176 => (( 5890.473, 4770.928),( 5875.455, 4796.938),( 5890.473, 4822.950),( 5875.455, 4848.961),( 5875.455, 5048.998),( 5890.473, 5075.009),( 5875.455, 5101.020),( 5890.473, 5127.031)), -- tube 176
   177 => (( 5920.507, 4770.928),( 5905.490, 4796.938),( 5920.507, 4822.950),( 5905.490, 4848.961),( 5905.490, 5048.998),( 5920.507, 5075.009),( 5905.490, 5101.020),( 5920.507, 5127.031)), -- tube 177
   178 => (( 5950.542, 4770.928),( 5935.525, 4796.938),( 5950.542, 4822.950),( 5935.525, 4848.961),( 5935.525, 5048.998),( 5950.542, 5075.009),( 5935.525, 5101.020),( 5950.542, 5127.031)), -- tube 178
   179 => (( 5980.578, 4770.928),( 5965.560, 4796.938),( 5980.578, 4822.950),( 5965.560, 4848.961),( 5965.560, 5048.998),( 5980.578, 5075.009),( 5965.560, 5101.020),( 5980.578, 5127.031)), -- tube 179
   180 => (( 6010.612, 4770.928),( 5995.595, 4796.938),( 6010.612, 4822.950),( 5995.595, 4848.961),( 5995.595, 5048.998),( 6010.612, 5075.009),( 5995.595, 5101.020),( 6010.612, 5127.031)), -- tube 180
   181 => (( 6040.647, 4770.928),( 6025.630, 4796.938),( 6040.647, 4822.950),( 6025.630, 4848.961),( 6025.630, 5048.998),( 6040.647, 5075.009),( 6025.630, 5101.020),( 6040.647, 5127.031)), -- tube 181
   182 => (( 6070.683, 4770.928),( 6055.665, 4796.938),( 6070.683, 4822.950),( 6055.665, 4848.961),( 6055.665, 5048.998),( 6070.683, 5075.009),( 6055.665, 5101.020),( 6070.683, 5127.031)), -- tube 182
   183 => (( 6100.717, 4770.928),( 6085.700, 4796.938),( 6100.717, 4822.950),( 6085.700, 4848.961),( 6085.700, 5048.998),( 6100.717, 5075.009),( 6085.700, 5101.020),( 6100.717, 5127.031)), -- tube 183
   184 => (( 6130.752, 4770.928),( 6115.735, 4796.938),( 6130.752, 4822.950),( 6115.735, 4848.961),( 6115.735, 5048.998),( 6130.752, 5075.009),( 6115.735, 5101.020),( 6130.752, 5127.031)), -- tube 184
   185 => (( 6160.788, 4770.928),( 6145.770, 4796.938),( 6160.788, 4822.950),( 6145.770, 4848.961),( 6145.770, 5048.998),( 6160.788, 5075.009),( 6145.770, 5101.020),( 6160.788, 5127.031)), -- tube 185
   186 => (( 6190.822, 4770.928),( 6175.805, 4796.938),( 6190.822, 4822.950),( 6175.805, 4848.961),( 6175.805, 5048.998),( 6190.822, 5075.009),( 6175.805, 5101.020),( 6190.822, 5127.031)), -- tube 186
   187 => (( 6220.857, 4770.928),( 6205.840, 4796.938),( 6220.857, 4822.950),( 6205.840, 4848.961),( 6205.840, 5048.998),( 6220.857, 5075.009),( 6205.840, 5101.020),( 6220.857, 5127.031)), -- tube 187
   188 => (( 6250.893, 4770.928),( 6235.875, 4796.938),( 6250.893, 4822.950),( 6235.875, 4848.961),( 6235.875, 5048.998),( 6250.893, 5075.009),( 6235.875, 5101.020),( 6250.893, 5127.031)), -- tube 188
   189 => (( 6280.928, 4770.928),( 6265.910, 4796.938),( 6280.928, 4822.950),( 6265.910, 4848.961),( 6265.910, 5048.998),( 6280.928, 5075.009),( 6265.910, 5101.020),( 6280.928, 5127.031)), -- tube 189
   190 => (( 6310.962, 4770.928),( 6295.945, 4796.938),( 6310.962, 4822.950),( 6295.945, 4848.961),( 6295.945, 5048.998),( 6310.962, 5075.009),( 6295.945, 5101.020),( 6310.962, 5127.031)), -- tube 190
   191 => (( 6340.998, 4770.928),( 6325.980, 4796.938),( 6340.998, 4822.950),( 6325.980, 4848.961),( 6325.980, 5048.998),( 6340.998, 5075.009),( 6325.980, 5101.020),( 6340.998, 5127.031)), -- tube 191
   192 => (( 6371.033, 4770.928),( 6356.015, 4796.938),( 6371.033, 4822.950),( 6356.015, 4848.961),( 6356.015, 5048.998),( 6371.033, 5075.009),( 6356.015, 5101.020),( 6371.033, 5127.031)), -- tube 192
   193 => (( 6401.067, 4770.928),( 6386.050, 4796.938),( 6401.067, 4822.950),( 6386.050, 4848.961),( 6386.050, 5048.998),( 6401.067, 5075.009),( 6386.050, 5101.020),( 6401.067, 5127.031)), -- tube 193
   194 => (( 6431.103, 4770.928),( 6416.085, 4796.938),( 6431.103, 4822.950),( 6416.085, 4848.961),( 6416.085, 5048.998),( 6431.103, 5075.009),( 6416.085, 5101.020),( 6431.103, 5127.031)), -- tube 194
   195 => (( 6461.138, 4770.928),( 6446.120, 4796.938),( 6461.138, 4822.950),( 6446.120, 4848.961),( 6446.120, 5048.998),( 6461.138, 5075.009),( 6446.120, 5101.020),( 6461.138, 5127.031)), -- tube 195
   196 => (( 6491.172, 4770.928),( 6476.155, 4796.938),( 6491.172, 4822.950),( 6476.155, 4848.961),( 6476.155, 5048.998),( 6491.172, 5075.009),( 6476.155, 5101.020),( 6491.172, 5127.031)), -- tube 196
   197 => (( 6521.208, 4770.928),( 6506.190, 4796.938),( 6521.208, 4822.950),( 6506.190, 4848.961),( 6506.190, 5048.998),( 6521.208, 5075.009),( 6506.190, 5101.020),( 6521.208, 5127.031))  -- tube 197
  );
  constant tube_coordinates_mid :  tube_coord_side_aat (0 to MAX_TUBES_MID - 1)(0 to 5):= (
    --     layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       ,
     0 => ((  135.000, 6913.458),(  150.018, 6939.468),(  135.000, 6965.479),(  135.000, 7312.517),(  150.018, 7338.528),(  135.000, 7364.540)), -- tube   0
     1 => ((  165.000, 6913.458),(  180.018, 6939.468),(  165.000, 6965.479),(  165.000, 7312.517),(  180.018, 7338.528),(  165.000, 7364.540)), -- tube   1
     2 => ((  195.035, 6913.458),(  210.053, 6939.468),(  195.035, 6965.479),(  195.035, 7312.517),(  210.053, 7338.528),(  195.035, 7364.540)), -- tube   2
     3 => ((  225.070, 6913.458),(  240.087, 6939.468),(  225.070, 6965.479),(  225.070, 7312.517),(  240.087, 7338.528),(  225.070, 7364.540)), -- tube   3
     4 => ((  255.105, 6913.458),(  270.122, 6939.468),(  255.105, 6965.479),(  255.105, 7312.517),(  270.122, 7338.528),(  255.105, 7364.540)), -- tube   4
     5 => ((  285.140, 6913.458),(  300.158, 6939.468),(  285.140, 6965.479),(  285.140, 7312.517),(  300.158, 7338.528),(  285.140, 7364.540)), -- tube   5
     6 => ((  315.175, 6913.458),(  330.193, 6939.468),(  315.175, 6965.479),(  315.175, 7312.517),(  330.193, 7338.528),(  315.175, 7364.540)), -- tube   6
     7 => ((  345.210, 6913.458),(  360.228, 6939.468),(  345.210, 6965.479),(  345.210, 7312.517),(  360.228, 7338.528),(  345.210, 7364.540)), -- tube   7
     8 => ((  375.245, 6913.458),(  390.263, 6939.468),(  375.245, 6965.479),(  375.245, 7312.517),(  390.263, 7338.528),(  375.245, 7364.540)), -- tube   8
     9 => ((  405.280, 6913.458),(  420.297, 6939.468),(  405.280, 6965.479),(  405.280, 7312.517),(  420.297, 7338.528),(  405.280, 7364.540)), -- tube   9
    10 => ((  435.315, 6913.458),(  450.332, 6939.468),(  435.315, 6965.479),(  435.315, 7312.517),(  450.332, 7338.528),(  435.315, 7364.540)), -- tube  10
    11 => ((  465.350, 6913.458),(  480.367, 6939.468),(  465.350, 6965.479),(  465.350, 7312.517),(  480.367, 7338.528),(  465.350, 7364.540)), -- tube  11
    12 => ((  495.385, 6913.458),(  510.402, 6939.468),(  495.385, 6965.479),(  495.385, 7312.517),(  510.402, 7338.528),(  495.385, 7364.540)), -- tube  12
    13 => ((  525.420, 6913.458),(  540.438, 6939.468),(  525.420, 6965.479),(  525.455, 7312.517),(  540.438, 7338.528),(  525.420, 7364.540)), -- tube  13
    14 => ((  555.455, 6913.458),(  570.472, 6939.468),(  555.455, 6965.479),(  555.455, 7312.517),(  570.472, 7338.528),(  555.455, 7364.540)), -- tube  14
    15 => ((  585.525, 6913.458),(  600.508, 6939.468),(  585.490, 6965.479),(  585.525, 7312.517),(  600.508, 7338.528),(  585.490, 7364.540)), -- tube  15
    16 => ((  615.525, 6913.458),(  630.542, 6939.468),(  615.525, 6965.479),(  615.525, 7312.517),(  630.542, 7338.528),(  615.525, 7364.540)), -- tube  16
    17 => ((  645.560, 6913.458),(  660.578, 6939.468),(  645.560, 6965.479),(  645.560, 7312.517),(  660.578, 7338.528),(  645.560, 7364.540)), -- tube  17
    18 => ((  675.595, 6913.458),(  690.612, 6939.468),(  675.595, 6965.479),(  675.595, 7312.517),(  690.612, 7338.528),(  675.595, 7364.540)), -- tube  18
    19 => ((  705.630, 6913.458),(  720.648, 6939.468),(  705.630, 6965.479),(  705.630, 7312.517),(  720.648, 7338.528),(  705.630, 7364.540)), -- tube  19
    20 => ((  735.665, 6913.458),(  750.682, 6939.468),(  735.665, 6965.479),(  735.665, 7312.517),(  750.682, 7338.528),(  735.665, 7364.540)), -- tube  20
    21 => ((  765.700, 6913.458),(  780.717, 6939.468),(  765.700, 6965.479),(  765.700, 7312.517),(  780.717, 7338.528),(  765.700, 7364.540)), -- tube  21
    22 => ((  795.735, 6913.458),(  810.753, 6939.468),(  795.735, 6965.479),(  795.735, 7312.517),(  810.753, 7338.528),(  795.735, 7364.540)), -- tube  22
    23 => ((  825.770, 6913.458),(  840.787, 6939.468),(  825.770, 6965.479),(  825.770, 7312.517),(  840.787, 7338.528),(  825.770, 7364.540)), -- tube  23
    24 => ((  855.805, 6913.458),(  870.823, 6939.468),(  855.805, 6965.479),(  855.805, 7312.517),(  870.857, 7338.528),(  855.805, 7364.540)), -- tube  24
    25 => ((  885.840, 6913.458),(  900.857, 6939.468),(  885.840, 6965.479),(  885.840, 7312.517),(  900.857, 7338.528),(  885.840, 7364.540)), -- tube  25
    26 => ((  915.875, 6913.458),(  930.893, 6939.468),(  915.875, 6965.479),(  915.875, 7312.517),(  930.857, 7338.528),(  915.875, 7364.540)), -- tube  26
    27 => ((  945.910, 6913.458),(  960.927, 6939.468),(  945.910, 6965.479),(  945.910, 7312.517),(  960.963, 7338.528),(  945.910, 7364.540)), -- tube  27
    28 => ((  975.945, 6913.458),(  990.963, 6939.468),(  975.945, 6965.479),(  975.980, 7312.517),(  990.963, 7338.528),(  975.945, 7364.540)), -- tube  28
    29 => (( 1006.015, 6913.458),( 1020.997, 6939.468),( 1005.980, 6965.479),( 1005.980, 7312.517),( 1020.997, 7338.528),( 1005.980, 7364.540)), -- tube  29
    30 => (( 1036.015, 6913.458),( 1051.032, 6939.468),( 1036.015, 6965.479),( 1036.015, 7312.517),( 1051.032, 7338.528),( 1036.015, 7364.540)), -- tube  30
    31 => (( 1066.050, 6913.458),( 1081.068, 6939.468),( 1066.050, 6965.479),( 1066.050, 7312.517),( 1081.068, 7338.528),( 1066.050, 7364.540)), -- tube  31
    32 => (( 1096.085, 6913.458),( 1111.103, 6939.468),( 1096.085, 6965.479),( 1096.085, 7312.517),( 1111.103, 7338.528),( 1096.085, 7364.540)), -- tube  32
    33 => (( 1126.120, 6913.458),( 1141.137, 6939.468),( 1126.120, 6965.479),( 1126.120, 7312.517),( 1141.137, 7338.528),( 1126.120, 7364.540)), -- tube  33
    34 => (( 1156.155, 6913.458),( 1171.172, 6939.468),( 1156.155, 6965.479),( 1156.155, 7312.517),( 1171.172, 7338.528),( 1156.155, 7364.540)), -- tube  34
    35 => (( 1186.190, 6913.458),( 1201.208, 6939.468),( 1186.190, 6965.479),( 1186.190, 7312.517),( 1201.208, 7338.528),( 1186.190, 7364.540)), -- tube  35
    36 => (( 1216.225, 6913.458),( 1231.243, 6939.468),( 1216.225, 6965.479),( 1216.225, 7312.517),( 1231.243, 7338.528),( 1216.225, 7364.540)), -- tube  36
    37 => (( 1246.260, 6913.458),( 1261.277, 6939.468),( 1246.260, 6965.479),( 1246.295, 7312.517),( 1261.277, 7338.528),( 1246.260, 7364.540)), -- tube  37
    38 => (( 1276.295, 6913.458),( 1291.312, 6939.468),( 1276.295, 6965.479),( 1276.295, 7312.517),( 1291.312, 7338.528),( 1276.295, 7364.540)), -- tube  38
    39 => (( 1306.330, 6913.458),( 1321.348, 6939.468),( 1306.330, 6965.479),( 1306.330, 7312.517),( 1321.348, 7338.528),( 1306.330, 7364.540)), -- tube  39
    40 => (( 1336.365, 6913.458),( 1351.382, 6939.468),( 1336.365, 6965.479),( 1336.365, 7312.517),( 1351.382, 7338.528),( 1336.365, 7364.540)), -- tube  40
    41 => (( 1366.400, 6913.458),( 1381.417, 6939.468),( 1366.400, 6965.479),( 1366.400, 7312.517),( 1381.417, 7338.528),( 1366.400, 7364.540)), -- tube  41
    42 => (( 1396.435, 6913.458),( 1411.453, 6939.468),( 1396.435, 6965.479),( 1396.435, 7312.517),( 1411.453, 7338.528),( 1396.435, 7364.540)), -- tube  42
    43 => (( 1426.470, 6913.458),( 1441.488, 6939.468),( 1426.470, 6965.479),( 1426.470, 7312.517),( 1441.488, 7338.528),( 1426.470, 7364.540)), -- tube  43
    44 => (( 1456.505, 6913.458),( 1471.522, 6939.468),( 1456.505, 6965.479),( 1456.505, 7312.517),( 1471.522, 7338.528),( 1456.505, 7364.540)), -- tube  44
    45 => (( 1486.540, 6913.458),( 1501.557, 6939.468),( 1486.540, 6965.479),( 1486.540, 7312.517),( 1501.557, 7338.528),( 1486.540, 7364.540)), -- tube  45
    46 => (( 1516.575, 6913.458),( 1531.593, 6939.468),( 1516.575, 6965.479),( 1516.575, 7312.517),( 1531.627, 7338.528),( 1516.575, 7364.540)), -- tube  46
    47 => (( 1546.610, 6913.458),( 1561.627, 6939.468),( 1546.610, 6965.479),( 1546.645, 7312.517),( 1561.627, 7338.528),( 1546.610, 7364.540)), -- tube  47
    48 => (( 1576.645, 6913.458),( 1591.662, 6939.468),( 1576.645, 6965.479),( 1576.645, 7312.517),( 1591.662, 7338.528),( 1576.645, 7364.540)), -- tube  48
    49 => (( 1606.680, 6913.458),( 1621.698, 6939.468),( 1606.680, 6965.479),( 1606.680, 7312.517),( 1621.698, 7338.528),( 1606.680, 7364.540)), -- tube  49
    50 => (( 1636.715, 6913.458),( 1651.733, 6939.468),( 1636.715, 6965.479),( 1636.750, 7312.517),( 1651.733, 7338.528),( 1636.715, 7364.540)), -- tube  50
    51 => (( 1666.750, 6913.458),( 1681.767, 6939.468),( 1666.750, 6965.479),( 1666.750, 7312.517),( 1681.767, 7338.528),( 1666.785, 7364.540)), -- tube  51
    52 => (( 1696.785, 6913.458),( 1711.802, 6939.468),( 1696.785, 6965.479),( 1696.785, 7312.517),( 1711.802, 7338.528),( 1696.785, 7364.540)), -- tube  52
    53 => (( 1726.820, 6913.458),( 1741.838, 6939.468),( 1726.820, 6965.479),( 1726.820, 7312.517),( 1741.838, 7338.528),( 1726.820, 7364.540)), -- tube  53
    54 => (( 1756.855, 6913.458),( 1771.872, 6939.468),( 1756.855, 6965.479),( 1756.855, 7312.517),( 1771.872, 7338.528),( 1756.855, 7364.540)), -- tube  54
    55 => (( 1786.890, 6913.458),( 1801.907, 6939.468),( 1786.890, 6965.479),( 1786.890, 7312.517),( 1801.907, 7338.528),( 1786.890, 7364.540)), -- tube  55
    56 => (( 1816.925, 6913.458),( 1831.943, 6939.468),( 1816.925, 6965.479),( 1816.925, 7312.517),( 1831.943, 7338.528),( 1816.925, 7364.540)), -- tube  56
    57 => (( 1865.000, 6913.458),( 1880.017, 6939.468),( 1865.000, 6965.479),( 1865.000, 7312.517),( 1880.017, 7338.528),( 1865.035, 7364.540)), -- tube  57
    58 => (( 1895.035, 6913.458),( 1910.052, 6939.468),( 1895.035, 6965.479),( 1895.035, 7312.517),( 1910.052, 7338.528),( 1895.035, 7364.540)), -- tube  58
    59 => (( 1925.070, 6913.458),( 1940.088, 6939.468),( 1925.070, 6965.479),( 1925.070, 7312.517),( 1940.088, 7338.528),( 1925.070, 7364.540)), -- tube  59
    60 => (( 1955.105, 6913.458),( 1970.123, 6939.468),( 1955.105, 6965.479),( 1955.105, 7312.517),( 1970.123, 7338.528),( 1955.105, 7364.540)), -- tube  60
    61 => (( 1985.140, 6913.458),( 2000.157, 6939.468),( 1985.140, 6965.479),( 1985.140, 7312.517),( 2000.157, 7338.528),( 1985.140, 7364.540)), -- tube  61
    62 => (( 2015.175, 6913.458),( 2030.193, 6939.468),( 2015.175, 6965.479),( 2015.175, 7312.517),( 2030.193, 7338.528),( 2015.210, 7364.540)), -- tube  62
    63 => (( 2045.210, 6913.458),( 2060.228, 6939.468),( 2045.210, 6965.479),( 2045.210, 7312.517),( 2060.228, 7338.528),( 2045.210, 7364.540)), -- tube  63
    64 => (( 2075.245, 6913.458),( 2090.262, 6939.468),( 2075.245, 6965.479),( 2075.245, 7312.517),( 2090.262, 7338.528),( 2075.245, 7364.540)), -- tube  64
    65 => (( 2105.280, 6913.458),( 2120.298, 6939.468),( 2105.280, 6965.479),( 2105.280, 7312.517),( 2120.298, 7338.528),( 2105.280, 7364.540)), -- tube  65
    66 => (( 2135.315, 6913.458),( 2150.333, 6939.468),( 2135.315, 6965.479),( 2135.315, 7312.517),( 2150.333, 7338.528),( 2135.315, 7364.540)), -- tube  66
    67 => (( 2165.350, 6913.458),( 2180.367, 6939.468),( 2165.350, 6965.479),( 2165.350, 7312.517),( 2180.367, 7338.528),( 2165.350, 7364.540)), -- tube  67
    68 => (( 2195.385, 6913.458),( 2210.403, 6939.468),( 2195.385, 6965.479),( 2195.385, 7312.517),( 2210.403, 7338.528),( 2195.385, 7364.540)), -- tube  68
    69 => (( 2225.420, 6913.458),( 2240.438, 6939.468),( 2225.420, 6965.479),( 2225.420, 7312.517),( 2240.438, 7338.528),( 2225.420, 7364.540)), -- tube  69
    70 => (( 2255.455, 6913.458),( 2270.472, 6939.468),( 2255.455, 6965.479),( 2255.455, 7312.517),( 2270.472, 7338.528),( 2255.455, 7364.540)), -- tube  70
    71 => (( 2285.490, 6913.458),( 2300.508, 6939.468),( 2285.490, 6965.479),( 2285.490, 7312.517),( 2300.508, 7338.528),( 2285.490, 7364.540)), -- tube  71
    72 => (( 2315.525, 6913.458),( 2330.542, 6939.468),( 2315.525, 6965.479),( 2315.525, 7312.517),( 2330.542, 7338.528),( 2315.525, 7364.540)), -- tube  72
    73 => (( 2345.560, 6913.458),( 2360.577, 6939.468),( 2345.560, 6965.479),( 2345.560, 7312.517),( 2360.577, 7338.528),( 2345.560, 7364.540)), -- tube  73
    74 => (( 2375.595, 6913.458),( 2390.613, 6939.468),( 2375.595, 6965.479),( 2375.595, 7312.517),( 2390.613, 7338.528),( 2375.595, 7364.540)), -- tube  74
    75 => (( 2405.630, 6913.458),( 2420.647, 6939.468),( 2405.630, 6965.479),( 2405.630, 7312.517),( 2420.647, 7338.528),( 2405.630, 7364.540)), -- tube  75
    76 => (( 2435.665, 6913.458),( 2450.683, 6939.468),( 2435.665, 6965.479),( 2435.665, 7312.517),( 2450.683, 7338.528),( 2435.665, 7364.540)), -- tube  76
    77 => (( 2465.700, 6913.458),( 2480.718, 6939.468),( 2465.700, 6965.479),( 2465.700, 7312.517),( 2480.718, 7338.528),( 2465.700, 7364.540)), -- tube  77
    78 => (( 2495.735, 6913.458),( 2510.752, 6939.468),( 2495.735, 6965.479),( 2495.735, 7312.517),( 2510.752, 7338.528),( 2495.735, 7364.540)), -- tube  78
    79 => (( 2525.770, 6913.458),( 2540.788, 6939.468),( 2525.770, 6965.479),( 2525.770, 7312.517),( 2540.788, 7338.528),( 2525.770, 7364.540)), -- tube  79
    80 => (( 2555.805, 6913.458),( 2570.823, 6939.468),( 2555.805, 6965.479),( 2555.805, 7312.517),( 2570.823, 7338.528),( 2555.805, 7364.540)), -- tube  80
    81 => (( 2585.840, 6913.458),( 2600.857, 6939.468),( 2585.840, 6965.479),( 2585.840, 7312.517),( 2600.857, 7338.528),( 2585.840, 7364.540)), -- tube  81
    82 => (( 2615.875, 6913.458),( 2630.893, 6939.468),( 2615.875, 6965.479),( 2615.875, 7312.517),( 2630.893, 7338.528),( 2615.875, 7364.540)), -- tube  82
    83 => (( 2645.910, 6913.458),( 2660.927, 6939.468),( 2645.910, 6965.479),( 2645.910, 7312.517),( 2660.927, 7338.528),( 2645.910, 7364.540)), -- tube  83
    84 => (( 2675.945, 6913.458),( 2690.962, 6939.468),( 2675.945, 6965.479),( 2675.945, 7312.517),( 2690.962, 7338.528),( 2675.945, 7364.540)), -- tube  84
    85 => (( 2705.980, 6913.458),( 2720.998, 6939.468),( 2705.980, 6965.479),( 2705.980, 7312.517),( 2720.998, 7338.528),( 2705.980, 7364.540)), -- tube  85
    86 => (( 2736.015, 6913.458),( 2751.032, 6939.468),( 2736.015, 6965.479),( 2736.015, 7312.517),( 2751.032, 7338.528),( 2736.015, 7364.540)), -- tube  86
    87 => (( 2766.050, 6913.458),( 2781.067, 6939.468),( 2766.050, 6965.479),( 2766.085, 7312.517),( 2781.067, 7338.528),( 2766.050, 7364.540)), -- tube  87
    88 => (( 2796.085, 6913.458),( 2811.103, 6939.468),( 2796.085, 6965.479),( 2796.085, 7312.517),( 2811.103, 7338.528),( 2796.085, 7364.540)), -- tube  88
    89 => (( 2826.120, 6913.458),( 2841.137, 6939.468),( 2826.120, 6965.479),( 2826.120, 7312.517),( 2841.137, 7338.528),( 2826.155, 7364.540)), -- tube  89
    90 => (( 2856.155, 6913.458),( 2871.173, 6939.468),( 2856.155, 6965.479),( 2856.155, 7312.517),( 2871.173, 7338.528),( 2856.155, 7364.540)), -- tube  90
    91 => (( 2886.190, 6913.458),( 2901.208, 6939.468),( 2886.190, 6965.479),( 2886.190, 7312.517),( 2901.208, 7338.528),( 2886.190, 7364.540)), -- tube  91
    92 => (( 2916.225, 6913.458),( 2931.242, 6939.468),( 2916.225, 6965.479),( 2916.225, 7312.517),( 2931.242, 7338.528),( 2916.225, 7364.540)), -- tube  92
    93 => (( 2946.260, 6913.458),( 2961.278, 6939.468),( 2946.260, 6965.479),( 2946.295, 7312.517),( 2961.278, 7338.528),( 2946.260, 7364.540)), -- tube  93
    94 => (( 2976.295, 6913.458),( 2991.312, 6939.468),( 2976.295, 6965.479),( 2976.295, 7312.517),( 2991.312, 7338.528),( 2976.295, 7364.540)), -- tube  94
    95 => (( 3006.330, 6913.458),( 3021.347, 6939.468),( 3006.330, 6965.479),( 3006.330, 7312.517),( 3021.347, 7338.528),( 3006.330, 7364.540)), -- tube  95
    96 => (( 3036.365, 6913.458),( 3051.383, 6939.468),( 3036.365, 6965.479),( 3036.365, 7312.517),( 3051.383, 7338.528),( 3036.365, 7364.540)), -- tube  96
    97 => (( 3066.400, 6913.458),( 3081.417, 6939.468),( 3066.400, 6965.479),( 3066.400, 7312.517),( 3081.417, 7338.528),( 3066.400, 7364.540)), -- tube  97
    98 => (( 3096.435, 6913.458),( 3111.452, 6939.468),( 3096.435, 6965.479),( 3096.435, 7312.517),( 3111.452, 7338.528),( 3096.435, 7364.540)), -- tube  98
    99 => (( 3126.470, 6913.458),( 3141.488, 6939.468),( 3126.470, 6965.479),( 3126.470, 7312.517),( 3141.488, 7338.528),( 3126.470, 7364.540)), -- tube  99
   100 => (( 3156.505, 6913.458),( 3171.522, 6939.468),( 3156.505, 6965.479),( 3156.505, 7312.517),( 3171.522, 7338.528),( 3156.505, 7364.540)), -- tube 100
   101 => (( 3186.540, 6913.458),( 3201.557, 6939.468),( 3186.540, 6965.479),( 3186.540, 7312.517),( 3201.557, 7338.528),( 3186.540, 7364.540)), -- tube 101
   102 => (( 3216.575, 6913.458),( 3231.593, 6939.468),( 3216.575, 6965.479),( 3216.575, 7312.517),( 3231.593, 7338.528),( 3216.575, 7364.540)), -- tube 102
   103 => (( 3246.610, 6913.458),( 3261.627, 6939.468),( 3246.610, 6965.479),( 3246.610, 7312.517),( 3261.627, 7338.528),( 3246.610, 7364.540)), -- tube 103
   104 => (( 3276.645, 6913.458),( 3291.663, 6939.468),( 3276.645, 6965.479),( 3276.645, 7312.517),( 3291.663, 7338.528),( 3276.645, 7364.540)), -- tube 104
   105 => (( 3306.680, 6913.458),( 3321.698, 6939.468),( 3306.680, 6965.479),( 3306.680, 7312.517),( 3321.698, 7338.528),( 3306.680, 7364.540)), -- tube 105
   106 => (( 3336.715, 6913.458),( 3351.732, 6939.468),( 3336.715, 6965.479),( 3336.715, 7312.517),( 3351.732, 7338.528),( 3336.715, 7364.540)), -- tube 106
   107 => (( 3366.750, 6913.458),( 3381.768, 6939.468),( 3366.750, 6965.479),( 3366.750, 7312.517),( 3381.768, 7338.528),( 3366.750, 7364.540)), -- tube 107
   108 => (( 3396.785, 6913.458),( 3411.802, 6939.468),( 3396.785, 6965.479),( 3396.785, 7312.517),( 3411.802, 7338.528),( 3396.785, 7364.540)), -- tube 108
   109 => (( 3426.820, 6913.458),( 3441.837, 6939.468),( 3426.820, 6965.479),( 3426.820, 7312.517),( 3441.837, 7338.528),( 3426.820, 7364.540)), -- tube 109
   110 => (( 3456.855, 6913.458),( 3471.873, 6939.468),( 3456.855, 6965.479),( 3456.855, 7312.517),( 3471.873, 7338.528),( 3456.855, 7364.540)), -- tube 110
   111 => (( 3486.890, 6913.458),( 3501.907, 6939.468),( 3486.890, 6965.479),( 3486.890, 7312.517),( 3501.907, 7338.528),( 3486.890, 7364.540)), -- tube 111
   112 => (( 3516.925, 6913.458),( 3531.942, 6939.468),( 3516.925, 6965.479),( 3516.925, 7312.517),( 3531.942, 7338.528),( 3516.925, 7364.540)), -- tube 112
   113 => (( 3565.000, 6913.458),( 3580.018, 6939.468),( 3565.000, 6965.479),( 3565.000, 7312.517),( 3580.018, 7338.528),( 3565.000, 7364.540)), -- tube 113
   114 => (( 3595.035, 6913.458),( 3610.052, 6939.468),( 3595.035, 6965.479),( 3595.035, 7312.517),( 3610.052, 7338.528),( 3595.035, 7364.540)), -- tube 114
   115 => (( 3625.070, 6913.458),( 3640.087, 6939.468),( 3625.070, 6965.479),( 3625.070, 7312.517),( 3640.087, 7338.528),( 3625.070, 7364.540)), -- tube 115
   116 => (( 3655.105, 6913.458),( 3670.123, 6939.468),( 3655.105, 6965.479),( 3655.105, 7312.517),( 3670.123, 7338.528),( 3655.105, 7364.540)), -- tube 116
   117 => (( 3685.140, 6913.458),( 3700.157, 6939.468),( 3685.140, 6965.479),( 3685.140, 7312.517),( 3700.157, 7338.528),( 3685.140, 7364.540)), -- tube 117
   118 => (( 3715.175, 6913.458),( 3730.192, 6939.468),( 3715.175, 6965.479),( 3715.175, 7312.517),( 3730.192, 7338.528),( 3715.175, 7364.540)), -- tube 118
   119 => (( 3745.210, 6913.458),( 3760.228, 6939.468),( 3745.210, 6965.479),( 3745.210, 7312.517),( 3760.228, 7338.528),( 3745.210, 7364.540)), -- tube 119
   120 => (( 3775.245, 6913.458),( 3790.262, 6939.468),( 3775.245, 6965.479),( 3775.245, 7312.517),( 3790.262, 7338.528),( 3775.245, 7364.540)), -- tube 120
   121 => (( 3805.280, 6913.458),( 3820.298, 6939.468),( 3805.280, 6965.479),( 3805.280, 7312.517),( 3820.298, 7338.528),( 3805.280, 7364.540)), -- tube 121
   122 => (( 3835.315, 6913.458),( 3850.333, 6939.468),( 3835.315, 6965.479),( 3835.315, 7312.517),( 3850.333, 7338.528),( 3835.315, 7364.540)), -- tube 122
   123 => (( 3865.350, 6913.458),( 3880.367, 6939.468),( 3865.350, 6965.479),( 3865.350, 7312.517),( 3880.367, 7338.528),( 3865.350, 7364.540)), -- tube 123
   124 => (( 3895.385, 6913.458),( 3910.403, 6939.468),( 3895.385, 6965.479),( 3895.385, 7312.517),( 3910.403, 7338.528),( 3895.385, 7364.540)), -- tube 124
   125 => (( 3925.420, 6913.458),( 3940.438, 6939.468),( 3925.420, 6965.479),( 3925.420, 7312.517),( 3940.438, 7338.528),( 3925.420, 7364.540)), -- tube 125
   126 => (( 3955.455, 6913.458),( 3970.472, 6939.468),( 3955.455, 6965.479),( 3955.455, 7312.517),( 3970.472, 7338.528),( 3955.455, 7364.540)), -- tube 126
   127 => (( 3985.490, 6913.458),( 4000.508, 6939.468),( 3985.490, 6965.479),( 3985.490, 7312.517),( 4000.508, 7338.528),( 3985.490, 7364.540)), -- tube 127
   128 => (( 4015.525, 6913.458),( 4030.542, 6939.468),( 4015.525, 6965.479),( 4015.525, 7312.517),( 4030.542, 7338.528),( 4015.525, 7364.540)), -- tube 128
   129 => (( 4045.560, 6913.458),( 4060.577, 6939.468),( 4045.560, 6965.479),( 4045.560, 7312.517),( 4060.577, 7338.528),( 4045.560, 7364.540)), -- tube 129
   130 => (( 4075.595, 6913.458),( 4090.613, 6939.468),( 4075.595, 6965.479),( 4075.595, 7312.517),( 4090.613, 7338.528),( 4075.595, 7364.540)), -- tube 130
   131 => (( 4105.630, 6913.458),( 4120.647, 6939.468),( 4105.630, 6965.479),( 4105.630, 7312.517),( 4120.647, 7338.528),( 4105.630, 7364.540)), -- tube 131
   132 => (( 4135.665, 6913.458),( 4150.683, 6939.468),( 4135.665, 6965.479),( 4135.665, 7312.517),( 4150.683, 7338.528),( 4135.665, 7364.540)), -- tube 132
   133 => (( 4165.700, 6913.458),( 4180.717, 6939.468),( 4165.700, 6965.479),( 4165.700, 7312.517),( 4180.717, 7338.528),( 4165.700, 7364.540)), -- tube 133
   134 => (( 4195.735, 6913.458),( 4210.752, 6939.468),( 4195.735, 6965.479),( 4195.735, 7312.517),( 4210.752, 7338.528),( 4195.735, 7364.540)), -- tube 134
   135 => (( 4225.770, 6913.458),( 4240.788, 6939.468),( 4225.770, 6965.479),( 4225.770, 7312.517),( 4240.788, 7338.528),( 4225.770, 7364.540)), -- tube 135
   136 => (( 4255.805, 6913.458),( 4270.822, 6939.468),( 4255.805, 6965.479),( 4255.805, 7312.517),( 4270.822, 7338.528),( 4255.805, 7364.540)), -- tube 136
   137 => (( 4285.840, 6913.458),( 4300.857, 6939.468),( 4285.840, 6965.479),( 4285.840, 7312.517),( 4300.857, 7338.528),( 4285.840, 7364.540)), -- tube 137
   138 => (( 4315.875, 6913.458),( 4330.893, 6939.468),( 4315.875, 6965.479),( 4315.875, 7312.517),( 4330.893, 7338.528),( 4315.875, 7364.540)), -- tube 138
   139 => (( 4345.910, 6913.458),( 4360.928, 6939.468),( 4345.910, 6965.479),( 4345.910, 7312.517),( 4360.928, 7338.528),( 4345.910, 7364.540)), -- tube 139
   140 => (( 4375.945, 6913.458),( 4390.962, 6939.468),( 4375.945, 6965.479),( 4375.945, 7312.517),( 4390.962, 7338.528),( 4375.945, 7364.540)), -- tube 140
   141 => (( 4405.980, 6913.458),( 4420.998, 6939.468),( 4405.980, 6965.479),( 4405.980, 7312.517),( 4420.998, 7338.528),( 4405.980, 7364.540)), -- tube 141
   142 => (( 4436.015, 6913.458),( 4451.033, 6939.468),( 4436.015, 6965.479),( 4436.015, 7312.517),( 4451.033, 7338.528),( 4436.015, 7364.540)), -- tube 142
   143 => (( 4466.050, 6913.458),( 4481.067, 6939.468),( 4466.050, 6965.479),( 4466.050, 7312.517),( 4481.067, 7338.528),( 4466.050, 7364.540)), -- tube 143
   144 => (( 4496.085, 6913.458),( 4511.103, 6939.468),( 4496.085, 6965.479),( 4496.085, 7312.517),( 4511.103, 7338.528),( 4496.085, 7364.540)), -- tube 144
   145 => (( 4526.120, 6913.458),( 4541.138, 6939.468),( 4526.120, 6965.479),( 4526.120, 7312.517),( 4541.138, 7338.528),( 4526.120, 7364.540)), -- tube 145
   146 => (( 4556.155, 6913.458),( 4571.172, 6939.468),( 4556.155, 6965.479),( 4556.155, 7312.517),( 4571.172, 7338.528),( 4556.155, 7364.540)), -- tube 146
   147 => (( 4586.190, 6913.458),( 4601.208, 6939.468),( 4586.190, 6965.479),( 4586.190, 7312.517),( 4601.208, 7338.528),( 4586.190, 7364.540)), -- tube 147
   148 => (( 4616.225, 6913.458),( 4631.243, 6939.468),( 4616.225, 6965.479),( 4616.225, 7312.517),( 4631.243, 7338.528),( 4616.225, 7364.540)), -- tube 148
   149 => (( 4646.260, 6913.458),( 4661.277, 6939.468),( 4646.260, 6965.479),( 4646.260, 7312.517),( 4661.277, 7338.528),( 4646.260, 7364.540)), -- tube 149
   150 => (( 4676.295, 6913.458),( 4691.312, 6939.468),( 4676.295, 6965.479),( 4676.295, 7312.517),( 4691.312, 7338.528),( 4676.295, 7364.540)), -- tube 150
   151 => (( 4706.330, 6913.458),( 4721.348, 6939.468),( 4706.330, 6965.479),( 4706.330, 7312.517),( 4721.348, 7338.528),( 4706.330, 7364.540)), -- tube 151
   152 => (( 4736.365, 6913.458),( 4751.382, 6939.468),( 4736.365, 6965.479),( 4736.365, 7312.517),( 4751.382, 7338.528),( 4736.365, 7364.540)), -- tube 152
   153 => (( 4766.400, 6913.458),( 4781.417, 6939.468),( 4766.400, 6965.479),( 4766.400, 7312.517),( 4781.417, 7338.528),( 4766.400, 7364.540)), -- tube 153
   154 => (( 4796.435, 6913.458),( 4811.453, 6939.468),( 4796.435, 6965.479),( 4796.435, 7312.517),( 4811.453, 7338.528),( 4796.435, 7364.540)), -- tube 154
   155 => (( 4826.470, 6913.458),( 4841.487, 6939.468),( 4826.470, 6965.479),( 4826.470, 7312.517),( 4841.487, 7338.528),( 4826.470, 7364.540)), -- tube 155
   156 => (( 4856.505, 6913.458),( 4871.522, 6939.468),( 4856.505, 6965.479),( 4856.505, 7312.517),( 4871.522, 7338.528),( 4856.505, 7364.540)), -- tube 156
   157 => (( 4886.540, 6913.458),( 4901.558, 6939.468),( 4886.540, 6965.479),( 4886.540, 7312.517),( 4901.558, 7338.528),( 4886.540, 7364.540)), -- tube 157
   158 => (( 4916.575, 6913.458),( 4931.592, 6939.468),( 4916.575, 6965.479),( 4916.575, 7312.517),( 4931.592, 7338.528),( 4916.575, 7364.540)), -- tube 158
   159 => (( 4946.610, 6913.458),( 4961.627, 6939.468),( 4946.610, 6965.479),( 4946.610, 7312.517),( 4961.627, 7338.528),( 4946.610, 7364.540)), -- tube 159
   160 => (( 4976.645, 6913.458),( 4991.663, 6939.468),( 4976.645, 6965.479),( 4976.645, 7312.517),( 4991.663, 7338.528),( 4976.645, 7364.540)), -- tube 160
   161 => (( 5006.680, 6913.458),( 5021.697, 6939.468),( 5006.680, 6965.479),( 5006.680, 7312.517),( 5021.697, 7338.528),( 5006.680, 7364.540)), -- tube 161
   162 => (( 5036.715, 6913.458),( 5051.732, 6939.468),( 5036.715, 6965.479),( 5036.715, 7312.517),( 5051.768, 7338.528),( 5036.715, 7364.540)), -- tube 162
   163 => (( 5066.750, 6913.458),( 5081.768, 6939.468),( 5066.750, 6965.479),( 5066.750, 7312.517),( 5081.768, 7338.528),( 5066.750, 7364.540)), -- tube 163
   164 => (( 5096.785, 6913.458),( 5111.803, 6939.468),( 5096.785, 6965.479),( 5096.785, 7312.517),( 5111.803, 7338.528),( 5096.785, 7364.540)), -- tube 164
   165 => (( 5126.820, 6913.458),( 5141.837, 6939.468),( 5126.820, 6965.479),( 5126.820, 7312.517),( 5141.837, 7338.528),( 5126.820, 7364.540)), -- tube 165
   166 => (( 5156.855, 6913.458),( 5171.873, 6939.468),( 5156.855, 6965.479),( 5156.855, 7312.517),( 5171.873, 7338.528),( 5156.855, 7364.540)), -- tube 166
   167 => (( 5186.890, 6913.458),( 5201.908, 6939.468),( 5186.890, 6965.479),( 5186.890, 7312.517),( 5201.908, 7338.528),( 5186.890, 7364.540)), -- tube 167
   168 => (( 5216.925, 6913.458),( 5231.942, 6939.468),( 5216.925, 6965.479),( 5216.925, 7312.517),( 5231.942, 7338.528),( 5216.925, 7364.540)), -- tube 168
   169 => (( 5265.000, 6913.458),( 5280.018, 6939.468),( 5265.000, 6965.479),( 5265.000, 7312.517),( 5280.018, 7338.528),( 5265.000, 7364.540)), -- tube 169
   170 => (( 5295.035, 6913.458),( 5310.053, 6939.468),( 5295.035, 6965.479),( 5295.035, 7312.517),( 5310.053, 7338.528),( 5295.035, 7364.540)), -- tube 170
   171 => (( 5325.070, 6913.458),( 5340.087, 6939.468),( 5325.070, 6965.479),( 5325.070, 7312.517),( 5340.087, 7338.528),( 5325.070, 7364.540)), -- tube 171
   172 => (( 5355.105, 6913.458),( 5370.123, 6939.468),( 5355.105, 6965.479),( 5355.105, 7312.517),( 5370.123, 7338.528),( 5355.105, 7364.540)), -- tube 172
   173 => (( 5385.140, 6913.458),( 5400.158, 6939.468),( 5385.140, 6965.479),( 5385.140, 7312.517),( 5400.158, 7338.528),( 5385.140, 7364.540)), -- tube 173
   174 => (( 5415.175, 6913.458),( 5430.192, 6939.468),( 5415.175, 6965.479),( 5415.175, 7312.517),( 5430.192, 7338.528),( 5415.175, 7364.540)), -- tube 174
   175 => (( 5445.210, 6913.458),( 5460.228, 6939.468),( 5445.210, 6965.479),( 5445.210, 7312.517),( 5460.228, 7338.528),( 5445.210, 7364.540)), -- tube 175
   176 => (( 5475.245, 6913.458),( 5490.263, 6939.468),( 5475.245, 6965.479),( 5475.245, 7312.517),( 5490.263, 7338.528),( 5475.245, 7364.540)), -- tube 176
   177 => (( 5505.280, 6913.458),( 5520.297, 6939.468),( 5505.280, 6965.479),( 5505.280, 7312.517),( 5520.297, 7338.528),( 5505.280, 7364.540)), -- tube 177
   178 => (( 5535.315, 6913.458),( 5550.333, 6939.468),( 5535.315, 6965.479),( 5535.315, 7312.517),( 5550.333, 7338.528),( 5535.315, 7364.540)), -- tube 178
   179 => (( 5565.350, 6913.458),( 5580.368, 6939.468),( 5565.350, 6965.479),( 5565.350, 7312.517),( 5580.368, 7338.528),( 5565.350, 7364.540)), -- tube 179
   180 => (( 5595.385, 6913.458),( 5610.402, 6939.468),( 5595.385, 6965.479),( 5595.385, 7312.517),( 5610.402, 7338.528),( 5595.385, 7364.540)), -- tube 180
   181 => (( 5625.420, 6913.458),( 5640.438, 6939.468),( 5625.420, 6965.479),( 5625.420, 7312.517),( 5640.438, 7338.528),( 5625.420, 7364.540)), -- tube 181
   182 => (( 5655.455, 6913.458),( 5670.473, 6939.468),( 5655.455, 6965.479),( 5655.455, 7312.517),( 5670.473, 7338.528),( 5655.455, 7364.540)), -- tube 182
   183 => (( 5685.490, 6913.458),( 5700.507, 6939.468),( 5685.490, 6965.479),( 5685.490, 7312.517),( 5700.507, 7338.528),( 5685.490, 7364.540)), -- tube 183
   184 => (( 5715.525, 6913.458),( 5730.542, 6939.468),( 5715.525, 6965.479),( 5715.525, 7312.517),( 5730.542, 7338.528),( 5715.525, 7364.540)), -- tube 184
   185 => (( 5745.560, 6913.458),( 5760.578, 6939.468),( 5745.560, 6965.479),( 5745.560, 7312.517),( 5760.578, 7338.528),( 5745.560, 7364.540)), -- tube 185
   186 => (( 5775.595, 6913.458),( 5790.612, 6939.468),( 5775.595, 6965.479),( 5775.595, 7312.517),( 5790.612, 7338.528),( 5775.595, 7364.540)), -- tube 186
   187 => (( 5805.630, 6913.458),( 5820.647, 6939.468),( 5805.630, 6965.479),( 5805.630, 7312.517),( 5820.647, 7338.528),( 5805.630, 7364.540)), -- tube 187
   188 => (( 5835.665, 6913.458),( 5850.683, 6939.468),( 5835.665, 6965.479),( 5835.665, 7312.517),( 5850.683, 7338.528),( 5835.665, 7364.540)), -- tube 188
   189 => (( 5865.700, 6913.458),( 5880.717, 6939.468),( 5865.700, 6965.479),( 5865.700, 7312.517),( 5880.717, 7338.528),( 5865.700, 7364.540)), -- tube 189
   190 => (( 5895.735, 6913.458),( 5910.752, 6939.468),( 5895.735, 6965.479),( 5895.735, 7312.517),( 5910.752, 7338.528),( 5895.735, 7364.540)), -- tube 190
   191 => (( 5925.770, 6913.458),( 5940.788, 6939.468),( 5925.770, 6965.479),( 5925.770, 7312.517),( 5940.788, 7338.528),( 5925.770, 7364.540)), -- tube 191
   192 => (( 5955.805, 6913.458),( 5970.822, 6939.468),( 5955.805, 6965.479),( 5955.805, 7312.517),( 5970.822, 7338.528),( 5955.805, 7364.540)), -- tube 192
   193 => (( 5985.840, 6913.458),( 6000.857, 6939.468),( 5985.840, 6965.479),( 5985.840, 7312.517),( 6000.857, 7338.528),( 5985.840, 7364.540)), -- tube 193
   194 => (( 6015.875, 6913.458),( 6030.893, 6939.468),( 6015.875, 6965.479),( 6015.875, 7312.517),( 6030.893, 7338.528),( 6015.875, 7364.540)), -- tube 194
   195 => (( 6045.910, 6913.458),( 6060.928, 6939.468),( 6045.910, 6965.479),( 6045.910, 7312.517),( 6060.928, 7338.528),( 6045.910, 7364.540)), -- tube 195
   196 => (( 6075.945, 6913.458),( 6090.962, 6939.468),( 6075.945, 6965.479),( 6075.945, 7312.517),( 6090.962, 7338.528),( 6075.945, 7364.540)), -- tube 196
   197 => (( 6105.980, 6913.458),( 6120.998, 6939.468),( 6105.980, 6965.479),( 6105.980, 7312.517),( 6120.998, 7338.528),( 6105.980, 7364.540)), -- tube 197
   198 => (( 6136.015, 6913.458),( 6151.033, 6939.468),( 6136.015, 6965.479),( 6136.015, 7312.517),( 6151.033, 7338.528),( 6136.015, 7364.540)), -- tube 198
   199 => (( 6166.050, 6913.458),( 6181.067, 6939.468),( 6166.050, 6965.479),( 6166.050, 7312.517),( 6181.067, 7338.528),( 6166.050, 7364.540)), -- tube 199
   200 => (( 6196.085, 6913.458),( 6211.103, 6939.468),( 6196.085, 6965.479),( 6196.085, 7312.517),( 6211.103, 7338.528),( 6196.085, 7364.540)), -- tube 200
   201 => (( 6226.120, 6913.458),( 6241.138, 6939.468),( 6226.120, 6965.479),( 6226.120, 7312.517),( 6241.138, 7338.528),( 6226.120, 7364.540)), -- tube 201
   202 => (( 6256.155, 6913.458),( 6271.172, 6939.468),( 6256.155, 6965.479),( 6256.155, 7312.517),( 6271.172, 7338.528),( 6256.155, 7364.540)), -- tube 202
   203 => (( 6286.190, 6913.458),( 6301.208, 6939.468),( 6286.190, 6965.479),( 6286.190, 7312.517),( 6301.208, 7338.528),( 6286.190, 7364.540)), -- tube 203
   204 => (( 6316.225, 6913.458),( 6331.243, 6939.468),( 6316.225, 6965.479),( 6316.225, 7312.517),( 6331.243, 7338.528),( 6316.225, 7364.540)), -- tube 204
   205 => (( 6346.260, 6913.458),( 6361.277, 6939.468),( 6346.260, 6965.479),( 6346.260, 7312.517),( 6361.277, 7338.528),( 6346.260, 7364.540)), -- tube 205
   206 => (( 6376.295, 6913.458),( 6391.312, 6939.468),( 6376.295, 6965.479),( 6376.295, 7312.517),( 6391.312, 7338.528),( 6376.295, 7364.540)), -- tube 206
   207 => (( 6406.330, 6913.458),( 6421.348, 6939.468),( 6406.330, 6965.479),( 6406.330, 7312.517),( 6421.348, 7338.528),( 6406.330, 7364.540)), -- tube 207
   208 => (( 6436.365, 6913.458),( 6451.382, 6939.468),( 6436.365, 6965.479),( 6436.365, 7312.517),( 6451.382, 7338.528),( 6436.365, 7364.540)), -- tube 208
   209 => (( 6485.000, 6913.458),( 6500.018, 6939.468),( 6485.000, 6965.479),( 6485.000, 7312.517),( 6500.018, 7338.528),( 6485.000, 7364.540)), -- tube 209
   210 => (( 6515.035, 6913.458),( 6530.053, 6939.468),( 6515.035, 6965.479),( 6515.035, 7312.517),( 6530.053, 7338.528),( 6515.035, 7364.540)), -- tube 210
   211 => (( 6545.070, 6913.458),( 6560.087, 6939.468),( 6545.070, 6965.479),( 6545.070, 7312.517),( 6560.087, 7338.528),( 6545.070, 7364.540)), -- tube 211
   212 => (( 6575.105, 6913.458),( 6590.123, 6939.468),( 6575.105, 6965.479),( 6575.105, 7312.517),( 6590.123, 7338.528),( 6575.105, 7364.540)), -- tube 212
   213 => (( 6605.140, 6913.458),( 6620.158, 6939.468),( 6605.140, 6965.479),( 6605.140, 7312.517),( 6620.158, 7338.528),( 6605.140, 7364.540)), -- tube 213
   214 => (( 6635.175, 6913.458),( 6650.192, 6939.468),( 6635.175, 6965.479),( 6635.175, 7312.517),( 6650.192, 7338.528),( 6635.175, 7364.540)), -- tube 214
   215 => (( 6665.210, 6913.458),( 6680.228, 6939.468),( 6665.210, 6965.479),( 6665.210, 7312.517),( 6680.228, 7338.528),( 6665.210, 7364.540)), -- tube 215
   216 => (( 6695.245, 6913.458),( 6710.263, 6939.468),( 6695.245, 6965.479),( 6695.245, 7312.517),( 6710.263, 7338.528),( 6695.245, 7364.540)), -- tube 216
   217 => (( 6725.280, 6913.458),( 6740.297, 6939.468),( 6725.280, 6965.479),( 6725.280, 7312.517),( 6740.297, 7338.528),( 6725.280, 7364.540)), -- tube 217
   218 => (( 6755.315, 6913.458),( 6770.333, 6939.468),( 6755.315, 6965.479),( 6755.315, 7312.517),( 6770.333, 7338.528),( 6755.315, 7364.540)), -- tube 218
   219 => (( 6785.350, 6913.458),( 6800.368, 6939.468),( 6785.350, 6965.479),( 6785.350, 7312.517),( 6800.368, 7338.528),( 6785.350, 7364.540)), -- tube 219
   220 => (( 6815.385, 6913.458),( 6830.402, 6939.468),( 6815.385, 6965.479),( 6815.385, 7312.517),( 6830.402, 7338.528),( 6815.385, 7364.540)), -- tube 220
   221 => (( 6845.420, 6913.458),( 6860.438, 6939.468),( 6845.420, 6965.479),( 6845.420, 7312.517),( 6860.438, 7338.528),( 6845.420, 7364.540)), -- tube 221
   222 => (( 6875.455, 6913.458),( 6890.473, 6939.468),( 6875.455, 6965.479),( 6875.455, 7312.517),( 6890.473, 7338.528),( 6875.455, 7364.540)), -- tube 222
   223 => (( 6905.490, 6913.458),( 6920.507, 6939.468),( 6905.490, 6965.479),( 6905.490, 7312.517),( 6920.507, 7338.528),( 6905.490, 7364.540)), -- tube 223
   224 => (( 6935.525, 6913.458),( 6950.542, 6939.468),( 6935.525, 6965.479),( 6935.525, 7312.517),( 6950.542, 7338.528),( 6935.525, 7364.540)), -- tube 224
   225 => (( 6965.560, 6913.458),( 6980.578, 6939.468),( 6965.560, 6965.479),( 6965.560, 7312.517),( 6980.578, 7338.528),( 6965.560, 7364.540)), -- tube 225
   226 => (( 6995.595, 6913.458),( 7010.612, 6939.468),( 6995.595, 6965.479),( 6995.595, 7312.517),( 7010.612, 7338.528),( 6995.595, 7364.540)), -- tube 226
   227 => (( 7025.630, 6913.458),( 7040.647, 6939.468),( 7025.630, 6965.479),( 7025.630, 7312.517),( 7040.647, 7338.528),( 7025.630, 7364.540)), -- tube 227
   228 => (( 7055.665, 6913.458),( 7070.683, 6939.468),( 7055.665, 6965.479),( 7055.665, 7312.517),( 7070.683, 7338.528),( 7055.665, 7364.540)), -- tube 228
   229 => (( 7085.700, 6913.458),( 7100.717, 6939.468),( 7085.700, 6965.479),( 7085.700, 7312.517),( 7100.717, 7338.528),( 7085.700, 7364.540)), -- tube 229
   230 => (( 7115.735, 6913.458),( 7130.752, 6939.468),( 7115.735, 6965.479),( 7115.735, 7312.517),( 7130.752, 7338.528),( 7115.735, 7364.540)), -- tube 230
   231 => (( 7145.770, 6913.458),( 7160.788, 6939.468),( 7145.770, 6965.479),( 7145.770, 7312.517),( 7160.788, 7338.528),( 7145.770, 7364.540)), -- tube 231
   232 => (( 7175.805, 6913.458),( 7190.822, 6939.468),( 7175.805, 6965.479),( 7175.805, 7312.517),( 7190.822, 7338.528),( 7175.805, 7364.540)), -- tube 232
   233 => (( 7205.840, 6913.458),( 7220.857, 6939.468),( 7205.840, 6965.479),( 7205.840, 7312.517),( 7220.857, 7338.528),( 7205.840, 7364.540)), -- tube 233
   234 => (( 7235.875, 6913.458),( 7250.893, 6939.468),( 7235.875, 6965.479),( 7235.875, 7312.517),( 7250.893, 7338.528),( 7235.875, 7364.540)), -- tube 234
   235 => (( 7265.910, 6913.458),( 7280.928, 6939.468),( 7265.910, 6965.479),( 7265.910, 7312.517),( 7280.928, 7338.528),( 7265.910, 7364.540)), -- tube 235
   236 => (( 7295.945, 6913.458),( 7310.962, 6939.468),( 7295.945, 6965.479),( 7295.945, 7312.517),( 7310.962, 7338.528),( 7295.945, 7364.540)), -- tube 236
   237 => (( 7325.980, 6913.458),( 7340.998, 6939.468),( 7325.980, 6965.479),( 7325.980, 7312.517),( 7340.998, 7338.528),( 7325.980, 7364.540)), -- tube 237
   238 => (( 7356.015, 6913.458),( 7371.033, 6939.468),( 7356.015, 6965.479),( 7356.015, 7312.517),( 7371.033, 7338.528),( 7356.015, 7364.540)), -- tube 238
   239 => (( 7386.050, 6913.458),( 7401.067, 6939.468),( 7386.050, 6965.479),( 7386.050, 7312.517),( 7401.067, 7338.528),( 7386.050, 7364.540)), -- tube 239
   240 => (( 7416.085, 6913.458),( 7431.103, 6939.468),( 7416.085, 6965.479),( 7416.085, 7312.517),( 7431.103, 7338.528),( 7416.085, 7364.540)), -- tube 240
   241 => (( 7446.120, 6913.458),( 7461.138, 6939.468),( 7446.120, 6965.479),( 7446.120, 7312.517),( 7461.138, 7338.528),( 7446.120, 7364.540)), -- tube 241
   242 => (( 7476.155, 6913.458),( 7491.172, 6939.468),( 7476.155, 6965.479),( 7476.155, 7312.517),( 7491.172, 7338.528),( 7476.155, 7364.540)), -- tube 242
   243 => (( 7506.190, 6913.458),( 7521.208, 6939.468),( 7506.190, 6965.479),( 7506.190, 7312.517),( 7521.208, 7338.528),( 7506.190, 7364.540)), -- tube 243
   244 => (( 7536.225, 6913.458),( 7551.243, 6939.468),( 7536.225, 6965.479),( 7536.225, 7312.517),( 7551.243, 7338.528),( 7536.225, 7364.540)), -- tube 244
   245 => (( 7566.260, 6913.458),( 7581.277, 6939.468),( 7566.260, 6965.479),( 7566.260, 7312.517),( 7581.277, 7338.528),( 7566.260, 7364.540)), -- tube 245
   246 => (( 7596.295, 6913.458),( 7611.312, 6939.468),( 7596.295, 6965.479),( 7596.295, 7312.517),( 7611.312, 7338.528),( 7596.295, 7364.540)), -- tube 246
   247 => (( 7626.330, 6913.458),( 7641.348, 6939.468),( 7626.330, 6965.479),( 7626.330, 7312.517),( 7641.348, 7338.528),( 7626.330, 7364.540)), -- tube 247
   248 => (( 7656.365, 6913.458),( 7671.382, 6939.468),( 7656.365, 6965.479),( 7656.365, 7312.517),( 7671.382, 7338.528),( 7656.365, 7364.540)), -- tube 248
   249 => (( 7705.000, 6913.458),( 7720.018, 6939.468),( 7705.000, 6965.479),( 7705.000, 7312.517),( 7720.018, 7338.528),( 7705.000, 7364.540)), -- tube 249
   250 => (( 7735.035, 6913.458),( 7750.053, 6939.468),( 7735.035, 6965.479),( 7735.035, 7312.517),( 7750.053, 7338.528),( 7735.035, 7364.540)), -- tube 250
   251 => (( 7765.070, 6913.458),( 7780.087, 6939.468),( 7765.070, 6965.479),( 7765.070, 7312.517),( 7780.087, 7338.528),( 7765.070, 7364.540)), -- tube 251
   252 => (( 7795.105, 6913.458),( 7810.123, 6939.468),( 7795.105, 6965.479),( 7795.105, 7312.517),( 7810.123, 7338.528),( 7795.105, 7364.540)), -- tube 252
   253 => (( 7825.140, 6913.458),( 7840.158, 6939.468),( 7825.140, 6965.479),( 7825.140, 7312.517),( 7840.158, 7338.528),( 7825.140, 7364.540)), -- tube 253
   254 => (( 7855.175, 6913.458),( 7870.192, 6939.468),( 7855.175, 6965.479),( 7855.175, 7312.517),( 7870.192, 7338.528),( 7855.175, 7364.540)), -- tube 254
   255 => (( 7885.210, 6913.458),( 7900.228, 6939.468),( 7885.210, 6965.479),( 7885.210, 7312.517),( 7900.228, 7338.528),( 7885.210, 7364.540)), -- tube 255
   256 => (( 7915.245, 6913.458),( 7930.263, 6939.468),( 7915.245, 6965.479),( 7915.245, 7312.517),( 7930.263, 7338.528),( 7915.245, 7364.540)), -- tube 256
   257 => (( 7945.280, 6913.458),( 7960.297, 6939.468),( 7945.280, 6965.479),( 7945.280, 7312.517),( 7960.297, 7338.528),( 7945.280, 7364.540)), -- tube 257
   258 => (( 7975.315, 6913.458),( 7990.333, 6939.468),( 7975.315, 6965.479),( 7975.315, 7312.517),( 7990.333, 7338.528),( 7975.315, 7364.540)), -- tube 258
   259 => (( 8005.350, 6913.458),( 8020.368, 6939.468),( 8005.350, 6965.479),( 8005.350, 7312.517),( 8020.368, 7338.528),( 8005.350, 7364.540)), -- tube 259
   260 => (( 8035.385, 6913.458),( 8050.402, 6939.468),( 8035.385, 6965.479),( 8035.385, 7312.517),( 8050.402, 7338.528),( 8035.385, 7364.540)), -- tube 260
   261 => (( 8065.420, 6913.458),( 8080.438, 6939.468),( 8065.420, 6965.479),( 8065.420, 7312.517),( 8080.438, 7338.528),( 8065.420, 7364.540)), -- tube 261
   262 => (( 8095.455, 6913.458),( 8110.473, 6939.468),( 8095.455, 6965.479),( 8095.455, 7312.517),( 8110.473, 7338.528),( 8095.455, 7364.540)), -- tube 262
   263 => (( 8125.490, 6913.458),( 8140.507, 6939.468),( 8125.490, 6965.479),( 8125.490, 7312.517),( 8140.507, 7338.528),( 8125.490, 7364.540)), -- tube 263
   264 => (( 8155.525, 6913.458),( 8170.542, 6939.468),( 8155.525, 6965.479),( 8155.525, 7312.517),( 8170.542, 7338.528),( 8155.525, 7364.540)), -- tube 264
   265 => (( 8185.560, 6913.458),( 8200.577, 6939.468),( 8185.560, 6965.479),( 8185.560, 7312.517),( 8200.577, 7338.528),( 8185.560, 7364.540)), -- tube 265
   266 => (( 8215.595, 6913.458),( 8230.612, 6939.468),( 8215.595, 6965.479),( 8215.595, 7312.517),( 8230.612, 7338.528),( 8215.595, 7364.540)), -- tube 266
   267 => (( 8245.630, 6913.458),( 8260.647, 6939.468),( 8245.630, 6965.479),( 8245.630, 7312.517),( 8260.647, 7338.528),( 8245.630, 7364.540)), -- tube 267
   268 => (( 8275.665, 6913.458),( 8290.683, 6939.468),( 8275.665, 6965.479),( 8275.665, 7312.517),( 8290.683, 7338.528),( 8275.665, 7364.540)), -- tube 268
   269 => (( 8305.700, 6913.458),( 8320.718, 6939.468),( 8305.700, 6965.479),( 8305.700, 7312.517),( 8320.718, 7338.528),( 8305.700, 7364.540)), -- tube 269
   270 => (( 8335.735, 6913.458),( 8350.753, 6939.468),( 8335.735, 6965.479),( 8335.735, 7312.517),( 8350.753, 7338.528),( 8335.735, 7364.540)), -- tube 270
   271 => (( 8365.770, 6913.458),( 8380.787, 6939.468),( 8365.770, 6965.479),( 8365.770, 7312.517),( 8380.787, 7338.528),( 8365.770, 7364.540)), -- tube 271
   272 => (( 8395.805, 6913.458),( 8410.822, 6939.468),( 8395.805, 6965.479),( 8395.805, 7312.517),( 8410.822, 7338.528),( 8395.805, 7364.540)), -- tube 272
   273 => (( 8425.840, 6913.458),( 8440.857, 6939.468),( 8425.840, 6965.479),( 8425.840, 7312.517),( 8440.857, 7338.528),( 8425.840, 7364.540)), -- tube 273
   274 => (( 8455.875, 6913.458),( 8470.893, 6939.468),( 8455.875, 6965.479),( 8455.875, 7312.517),( 8470.893, 7338.528),( 8455.875, 7364.540)), -- tube 274
   275 => (( 8485.910, 6913.458),( 8500.928, 6939.468),( 8485.910, 6965.479),( 8485.910, 7312.517),( 8500.928, 7338.528),( 8485.910, 7364.540)), -- tube 275
   276 => (( 8515.945, 6913.458),( 8530.963, 6939.468),( 8515.945, 6965.479),( 8515.945, 7312.517),( 8530.963, 7338.528),( 8515.945, 7364.540)), -- tube 276
   277 => (( 8545.980, 6913.458),( 8560.997, 6939.468),( 8545.980, 6965.479),( 8545.980, 7312.517),( 8560.997, 7338.528),( 8545.980, 7364.540)), -- tube 277
   278 => (( 8576.015, 6913.458),( 8591.032, 6939.468),( 8576.015, 6965.479),( 8576.015, 7312.517),( 8591.032, 7338.528),( 8576.015, 7364.540)), -- tube 278
   279 => (( 8606.050, 6913.458),( 8621.067, 6939.468),( 8606.050, 6965.479),( 8606.050, 7312.517),( 8621.067, 7338.528),( 8606.050, 7364.540)), -- tube 279
   280 => (( 8636.085, 6913.458),( 8651.103, 6939.468),( 8636.085, 6965.479),( 8636.085, 7312.517),( 8651.103, 7338.528),( 8636.085, 7364.540)), -- tube 280
   281 => (( 8666.120, 6913.458),( 8681.138, 6939.468),( 8666.120, 6965.479),( 8666.120, 7312.517),( 8681.138, 7338.528),( 8666.120, 7364.540)), -- tube 281
   282 => (( 8696.155, 6913.458),( 8711.173, 6939.468),( 8696.155, 6965.479),( 8696.155, 7312.517),( 8711.173, 7338.528),( 8696.155, 7364.540)), -- tube 282
   283 => (( 8726.190, 6913.458),( 8741.207, 6939.468),( 8726.190, 6965.479),( 8726.190, 7312.517),( 8741.207, 7338.528),( 8726.190, 7364.540)), -- tube 283
   284 => (( 8756.225, 6913.458),( 8771.242, 6939.468),( 8756.225, 6965.479),( 8756.225, 7312.517),( 8771.242, 7338.528),( 8756.225, 7364.540)), -- tube 284
   285 => (( 8786.260, 6913.458),( 8801.277, 6939.468),( 8786.260, 6965.479),( 8786.260, 7312.517),( 8801.277, 7338.528),( 8786.260, 7364.540)), -- tube 285
   286 => (( 8816.295, 6913.458),( 8831.312, 6939.468),( 8816.295, 6965.479),( 8816.295, 7312.517),( 8831.312, 7338.528),( 8816.295, 7364.540)), -- tube 286
   287 => (( 8846.330, 6913.458),( 8861.348, 6939.468),( 8846.330, 6965.479),( 8846.330, 7312.517),( 8861.348, 7338.528),( 8846.330, 7364.540)), -- tube 287
   288 => (( 8876.365, 6913.458),( 8891.383, 6939.468),( 8876.365, 6965.479),( 8876.365, 7312.517),( 8891.383, 7338.528),( 8876.365, 7364.540)), -- tube 288
   289 => (( 8906.400, 6913.458),( 8921.418, 6939.468),( 8906.400, 6965.479),( 8906.400, 7312.517),( 8921.418, 7338.528),( 8906.400, 7364.540)), -- tube 289
   290 => (( 8936.435, 6913.458),( 8951.452, 6939.468),( 8936.435, 6965.479),( 8936.435, 7312.517),( 8951.452, 7338.528),( 8936.435, 7364.540)), -- tube 290
   291 => (( 8966.470, 6913.458),( 8981.487, 6939.468),( 8966.470, 6965.479),( 8966.470, 7312.517),( 8981.487, 7338.528),( 8966.470, 7364.540)), -- tube 291
   292 => (( 8996.505, 6913.458),( 9011.522, 6939.468),( 8996.505, 6965.479),( 8996.505, 7312.517),( 9011.522, 7338.528),( 8996.505, 7364.540)), -- tube 292
   293 => (( 9026.540, 6913.458),( 9041.558, 6939.468),( 9026.540, 6965.479),( 9026.540, 7312.517),( 9041.558, 7338.528),( 9026.540, 7364.540)), -- tube 293
   294 => (( 9056.575, 6913.458),( 9071.593, 6939.468),( 9056.575, 6965.479),( 9056.575, 7312.517),( 9071.593, 7338.528),( 9056.575, 7364.540)), -- tube 294
   295 => (( 9086.610, 6913.458),( 9101.628, 6939.468),( 9086.610, 6965.479),( 9086.610, 7312.517),( 9101.628, 7338.528),( 9086.610, 7364.540))  -- tube 295
  );
  constant tube_coordinates_out :  tube_coord_side_aat (0 to MAX_TUBES_OUT - 1)(0 to 5):= (
    --      layer 0       , layer 1       , layer 2       , layer 3       , layer 4       , layer 5       ,
     0 => ((  135.000, 9274.457),(  150.018, 9300.469),(  135.000, 9326.479),(  135.000, 9673.518),(  150.018, 9699.528),(  135.000, 9725.539)), -- tube   0
     1 => ((  165.000, 9274.457),(  180.018, 9300.469),(  165.000, 9326.479),(  165.000, 9673.518),(  180.018, 9699.528),(  165.000, 9725.539)), -- tube   1
     2 => ((  195.035, 9274.457),(  210.053, 9300.469),(  195.035, 9326.479),(  195.035, 9673.518),(  210.087, 9699.528),(  195.035, 9725.539)), -- tube   2
     3 => ((  225.070, 9274.457),(  240.087, 9300.469),(  225.070, 9326.479),(  225.070, 9673.518),(  240.087, 9699.528),(  225.070, 9725.539)), -- tube   3
     4 => ((  255.105, 9274.457),(  270.122, 9300.469),(  255.105, 9326.479),(  255.105, 9673.518),(  270.122, 9699.528),(  255.105, 9725.539)), -- tube   4
     5 => ((  285.140, 9274.457),(  300.158, 9300.469),(  285.140, 9326.479),(  285.140, 9673.518),(  300.158, 9699.528),(  285.140, 9725.539)), -- tube   5
     6 => ((  315.175, 9274.457),(  330.193, 9300.469),(  315.175, 9326.479),(  315.175, 9673.518),(  330.193, 9699.528),(  315.175, 9725.539)), -- tube   6
     7 => ((  345.210, 9274.457),(  360.228, 9300.469),(  345.210, 9326.479),(  345.210, 9673.518),(  360.228, 9699.528),(  345.210, 9725.539)), -- tube   7
     8 => ((  375.245, 9274.457),(  390.263, 9300.469),(  375.245, 9326.479),(  375.245, 9673.518),(  390.263, 9699.528),(  375.245, 9725.539)), -- tube   8
     9 => ((  405.280, 9274.457),(  420.297, 9300.469),(  405.280, 9326.479),(  405.280, 9673.518),(  420.297, 9699.528),(  405.280, 9725.539)), -- tube   9
    10 => ((  435.315, 9274.457),(  450.332, 9300.469),(  435.315, 9326.479),(  435.350, 9673.518),(  450.332, 9699.528),(  435.315, 9725.539)), -- tube  10
    11 => ((  465.350, 9274.457),(  480.367, 9300.469),(  465.350, 9326.479),(  465.350, 9673.518),(  480.367, 9699.528),(  465.350, 9725.539)), -- tube  11
    12 => ((  495.385, 9274.457),(  510.402, 9300.469),(  495.385, 9326.479),(  495.385, 9673.518),(  510.402, 9699.528),(  495.385, 9725.539)), -- tube  12
    13 => ((  525.420, 9274.457),(  540.438, 9300.469),(  525.420, 9326.479),(  525.420, 9673.518),(  540.438, 9699.528),(  525.420, 9725.539)), -- tube  13
    14 => ((  555.455, 9274.457),(  570.472, 9300.469),(  555.455, 9326.479),(  555.455, 9673.518),(  570.472, 9699.528),(  555.490, 9725.539)), -- tube  14
    15 => ((  585.490, 9274.457),(  600.508, 9300.469),(  585.490, 9326.479),(  585.490, 9673.518),(  600.508, 9699.528),(  585.490, 9725.539)), -- tube  15
    16 => ((  615.525, 9274.457),(  630.542, 9300.469),(  615.525, 9326.479),(  615.525, 9673.518),(  630.542, 9699.528),(  615.525, 9725.539)), -- tube  16
    17 => ((  645.560, 9274.457),(  660.578, 9300.469),(  645.560, 9326.479),(  645.560, 9673.518),(  660.578, 9699.528),(  645.560, 9725.539)), -- tube  17
    18 => ((  675.595, 9274.457),(  690.612, 9300.469),(  675.595, 9326.479),(  675.595, 9673.518),(  690.612, 9699.528),(  675.630, 9725.539)), -- tube  18
    19 => ((  705.630, 9274.457),(  720.648, 9300.469),(  705.630, 9326.479),(  705.630, 9673.518),(  720.648, 9699.528),(  705.630, 9725.539)), -- tube  19
    20 => ((  735.665, 9274.457),(  750.682, 9300.469),(  735.665, 9326.479),(  735.665, 9673.518),(  750.682, 9699.528),(  735.665, 9725.539)), -- tube  20
    21 => ((  765.700, 9274.457),(  780.717, 9300.469),(  765.700, 9326.479),(  765.700, 9673.518),(  780.717, 9699.528),(  765.700, 9725.539)), -- tube  21
    22 => ((  795.735, 9274.457),(  810.753, 9300.469),(  795.735, 9326.479),(  795.735, 9673.518),(  810.753, 9699.528),(  795.735, 9725.539)), -- tube  22
    23 => ((  825.770, 9274.457),(  840.787, 9300.469),(  825.770, 9326.479),(  825.770, 9673.518),(  840.787, 9699.528),(  825.770, 9725.539)), -- tube  23
    24 => ((  855.805, 9274.457),(  870.823, 9300.469),(  855.805, 9326.479),(  855.805, 9673.518),(  870.823, 9699.528),(  855.805, 9725.539)), -- tube  24
    25 => ((  885.840, 9274.457),(  900.857, 9300.469),(  885.840, 9326.479),(  885.840, 9673.518),(  900.857, 9699.528),(  885.840, 9725.539)), -- tube  25
    26 => ((  915.875, 9274.457),(  930.893, 9300.469),(  915.875, 9326.479),(  915.875, 9673.518),(  930.893, 9699.528),(  915.875, 9725.539)), -- tube  26
    27 => ((  945.910, 9274.457),(  960.927, 9300.469),(  945.910, 9326.479),(  945.945, 9673.518),(  960.927, 9699.528),(  945.910, 9725.539)), -- tube  27
    28 => ((  975.945, 9274.457),(  990.963, 9300.469),(  975.945, 9326.479),(  975.945, 9673.518),(  990.963, 9699.528),(  975.945, 9725.539)), -- tube  28
    29 => (( 1005.980, 9274.457),( 1020.997, 9300.469),( 1005.980, 9326.479),( 1005.980, 9673.518),( 1020.997, 9699.528),( 1005.980, 9725.539)), -- tube  29
    30 => (( 1036.015, 9274.457),( 1051.032, 9300.469),( 1036.050, 9326.479),( 1036.015, 9673.518),( 1051.032, 9699.528),( 1036.015, 9725.539)), -- tube  30
    31 => (( 1066.050, 9274.457),( 1081.103, 9300.469),( 1066.050, 9326.479),( 1066.050, 9673.518),( 1081.068, 9699.528),( 1066.050, 9725.539)), -- tube  31
    32 => (( 1096.085, 9274.457),( 1111.103, 9300.469),( 1096.085, 9326.479),( 1096.085, 9673.518),( 1111.103, 9699.528),( 1096.085, 9725.539)), -- tube  32
    33 => (( 1126.120, 9274.457),( 1141.137, 9300.469),( 1126.120, 9326.479),( 1126.120, 9673.518),( 1141.137, 9699.528),( 1126.120, 9725.539)), -- tube  33
    34 => (( 1156.155, 9274.457),( 1171.172, 9300.469),( 1156.155, 9326.479),( 1156.155, 9673.518),( 1171.172, 9699.528),( 1156.155, 9725.539)), -- tube  34
    35 => (( 1186.225, 9274.457),( 1201.208, 9300.469),( 1186.190, 9326.479),( 1186.190, 9673.518),( 1201.208, 9699.528),( 1186.190, 9725.539)), -- tube  35
    36 => (( 1216.225, 9274.457),( 1231.243, 9300.469),( 1216.225, 9326.479),( 1216.225, 9673.518),( 1231.243, 9699.528),( 1216.225, 9725.539)), -- tube  36
    37 => (( 1246.260, 9274.457),( 1261.312, 9300.469),( 1246.260, 9326.479),( 1246.260, 9673.518),( 1261.277, 9699.528),( 1246.260, 9725.539)), -- tube  37
    38 => (( 1276.295, 9274.457),( 1291.312, 9300.469),( 1276.295, 9326.479),( 1276.295, 9673.518),( 1291.312, 9699.528),( 1276.295, 9725.539)), -- tube  38
    39 => (( 1306.330, 9274.457),( 1321.348, 9300.469),( 1306.330, 9326.479),( 1306.330, 9673.518),( 1321.348, 9699.528),( 1306.330, 9725.539)), -- tube  39
    40 => (( 1336.365, 9274.457),( 1351.382, 9300.469),( 1336.365, 9326.479),( 1336.365, 9673.518),( 1351.382, 9699.528),( 1336.365, 9725.539)), -- tube  40
    41 => (( 1366.400, 9274.457),( 1381.417, 9300.469),( 1366.400, 9326.479),( 1366.400, 9673.518),( 1381.417, 9699.528),( 1366.400, 9725.539)), -- tube  41
    42 => (( 1396.435, 9274.457),( 1411.453, 9300.469),( 1396.435, 9326.479),( 1396.435, 9673.518),( 1411.453, 9699.528),( 1396.435, 9725.539)), -- tube  42
    43 => (( 1426.470, 9274.457),( 1441.488, 9300.469),( 1426.470, 9326.479),( 1426.470, 9673.518),( 1441.488, 9699.528),( 1426.470, 9725.539)), -- tube  43
    44 => (( 1456.505, 9274.457),( 1471.522, 9300.469),( 1456.505, 9326.479),( 1456.505, 9673.518),( 1471.522, 9699.528),( 1456.505, 9725.539)), -- tube  44
    45 => (( 1486.540, 9274.457),( 1501.557, 9300.469),( 1486.540, 9326.479),( 1486.540, 9673.518),( 1501.557, 9699.528),( 1486.540, 9725.539)), -- tube  45
    46 => (( 1516.575, 9274.457),( 1531.593, 9300.469),( 1516.575, 9326.479),( 1516.575, 9673.518),( 1531.593, 9699.528),( 1516.575, 9725.539)), -- tube  46
    47 => (( 1546.610, 9274.457),( 1561.627, 9300.469),( 1546.610, 9326.479),( 1546.610, 9673.518),( 1561.627, 9699.528),( 1546.610, 9725.539)), -- tube  47
    48 => (( 1576.645, 9274.457),( 1591.662, 9300.469),( 1576.645, 9326.479),( 1576.645, 9673.518),( 1591.662, 9699.528),( 1576.645, 9725.539)), -- tube  48
    49 => (( 1606.680, 9274.457),( 1621.698, 9300.469),( 1606.680, 9326.479),( 1606.680, 9673.518),( 1621.698, 9699.528),( 1606.680, 9725.539)), -- tube  49
    50 => (( 1636.715, 9274.457),( 1651.733, 9300.469),( 1636.715, 9326.479),( 1636.715, 9673.518),( 1651.767, 9699.528),( 1636.715, 9725.539)), -- tube  50
    51 => (( 1666.750, 9274.457),( 1681.767, 9300.469),( 1666.750, 9326.479),( 1666.750, 9673.518),( 1681.767, 9699.528),( 1666.750, 9725.539)), -- tube  51
    52 => (( 1696.785, 9274.457),( 1711.802, 9300.469),( 1696.785, 9326.479),( 1696.785, 9673.518),( 1711.802, 9699.528),( 1696.785, 9725.539)), -- tube  52
    53 => (( 1726.820, 9274.457),( 1741.838, 9300.469),( 1726.820, 9326.479),( 1726.820, 9673.518),( 1741.838, 9699.528),( 1726.820, 9725.539)), -- tube  53
    54 => (( 1756.855, 9274.457),( 1771.872, 9300.469),( 1756.855, 9326.479),( 1756.855, 9673.518),( 1771.872, 9699.528),( 1756.855, 9725.539)), -- tube  54
    55 => (( 1786.890, 9274.457),( 1801.907, 9300.469),( 1786.890, 9326.479),( 1786.890, 9673.518),( 1801.943, 9699.528),( 1786.890, 9725.539)), -- tube  55
    56 => (( 1816.925, 9274.457),( 1831.943, 9300.469),( 1816.960, 9326.479),( 1816.925, 9673.518),( 1831.943, 9699.528),( 1816.925, 9725.539)), -- tube  56
    57 => (( 1846.960, 9274.457),( 1861.978, 9300.469),( 1846.960, 9326.479),( 1846.960, 9673.518),( 1861.978, 9699.528),( 1846.960, 9725.539)), -- tube  57
    58 => (( 1876.995, 9274.457),( 1892.012, 9300.469),( 1876.995, 9326.479),( 1876.995, 9673.518),( 1892.012, 9699.528),( 1876.995, 9725.539)), -- tube  58
    59 => (( 1907.030, 9274.457),( 1922.047, 9300.469),( 1907.030, 9326.479),( 1907.030, 9673.518),( 1922.047, 9699.528),( 1907.030, 9725.539)), -- tube  59
    60 => (( 1937.065, 9274.457),( 1952.083, 9300.469),( 1937.065, 9326.479),( 1937.065, 9673.518),( 1952.083, 9699.528),( 1937.065, 9725.539)), -- tube  60
    61 => (( 1967.100, 9274.457),( 1982.117, 9300.469),( 1967.100, 9326.479),( 1967.100, 9673.518),( 1982.117, 9699.528),( 1967.100, 9725.539)), -- tube  61
    62 => (( 1997.135, 9274.457),( 2012.152, 9300.469),( 1997.135, 9326.479),( 1997.135, 9673.518),( 2012.152, 9699.528),( 1997.135, 9725.539)), -- tube  62
    63 => (( 2027.170, 9274.457),( 2042.188, 9300.469),( 2027.170, 9326.479),( 2027.170, 9673.518),( 2042.188, 9699.528),( 2027.170, 9725.539)), -- tube  63
    64 => (( 2057.205, 9274.457),( 2072.222, 9300.469),( 2057.205, 9326.479),( 2057.205, 9673.518),( 2072.222, 9699.528),( 2057.205, 9725.539)), -- tube  64
    65 => (( 2087.240, 9274.457),( 2102.258, 9300.469),( 2087.240, 9326.479),( 2087.240, 9673.518),( 2102.258, 9699.528),( 2087.240, 9725.539)), -- tube  65
    66 => (( 2117.275, 9274.457),( 2132.292, 9300.469),( 2117.275, 9326.479),( 2117.275, 9673.518),( 2132.292, 9699.528),( 2117.275, 9725.539)), -- tube  66
    67 => (( 2147.310, 9274.457),( 2162.327, 9300.469),( 2147.310, 9326.479),( 2147.310, 9673.518),( 2162.327, 9699.528),( 2147.310, 9725.539)), -- tube  67
    68 => (( 2177.345, 9274.457),( 2192.363, 9300.469),( 2177.345, 9326.479),( 2177.345, 9673.518),( 2192.363, 9699.528),( 2177.345, 9725.539)), -- tube  68
    69 => (( 2207.380, 9274.457),( 2222.397, 9300.469),( 2207.380, 9326.479),( 2207.380, 9673.518),( 2222.397, 9699.528),( 2207.380, 9725.539)), -- tube  69
    70 => (( 2237.415, 9274.457),( 2252.432, 9300.469),( 2237.415, 9326.479),( 2237.415, 9673.518),( 2252.432, 9699.528),( 2237.415, 9725.539)), -- tube  70
    71 => (( 2267.450, 9274.457),( 2282.468, 9300.469),( 2267.450, 9326.479),( 2267.450, 9673.518),( 2282.468, 9699.528),( 2267.450, 9725.539)), -- tube  71
    72 => (( 2297.485, 9274.457),( 2312.502, 9300.469),( 2297.485, 9326.479),( 2297.485, 9673.518),( 2312.502, 9699.528),( 2297.485, 9725.539)), -- tube  72
    73 => (( 2345.000, 9274.457),( 2360.018, 9300.469),( 2345.000, 9326.479),( 2345.000, 9673.518),( 2360.018, 9699.528),( 2345.000, 9725.539)), -- tube  73
    74 => (( 2375.035, 9274.457),( 2390.052, 9300.469),( 2375.035, 9326.479),( 2375.035, 9673.518),( 2390.052, 9699.528),( 2375.035, 9725.539)), -- tube  74
    75 => (( 2405.070, 9274.457),( 2420.087, 9300.469),( 2405.070, 9326.479),( 2405.070, 9673.518),( 2420.087, 9699.528),( 2405.070, 9725.539)), -- tube  75
    76 => (( 2435.105, 9274.457),( 2450.123, 9300.469),( 2435.105, 9326.479),( 2435.105, 9673.518),( 2450.123, 9699.528),( 2435.105, 9725.539)), -- tube  76
    77 => (( 2465.140, 9274.457),( 2480.157, 9300.469),( 2465.140, 9326.479),( 2465.140, 9673.518),( 2480.157, 9699.528),( 2465.140, 9725.539)), -- tube  77
    78 => (( 2495.175, 9274.457),( 2510.192, 9300.469),( 2495.175, 9326.479),( 2495.175, 9673.518),( 2510.192, 9699.528),( 2495.175, 9725.539)), -- tube  78
    79 => (( 2525.210, 9274.457),( 2540.228, 9300.469),( 2525.210, 9326.479),( 2525.210, 9673.518),( 2540.228, 9699.528),( 2525.210, 9725.539)), -- tube  79
    80 => (( 2555.245, 9274.457),( 2570.262, 9300.469),( 2555.245, 9326.479),( 2555.245, 9673.518),( 2570.298, 9699.528),( 2555.245, 9725.539)), -- tube  80
    81 => (( 2585.280, 9274.457),( 2600.298, 9300.469),( 2585.280, 9326.479),( 2585.280, 9673.518),( 2600.298, 9699.528),( 2585.280, 9725.539)), -- tube  81
    82 => (( 2615.315, 9274.457),( 2630.333, 9300.469),( 2615.315, 9326.479),( 2615.315, 9673.518),( 2630.333, 9699.528),( 2615.315, 9725.539)), -- tube  82
    83 => (( 2645.350, 9274.457),( 2660.367, 9300.469),( 2645.350, 9326.479),( 2645.350, 9673.518),( 2660.367, 9699.528),( 2645.350, 9725.539)), -- tube  83
    84 => (( 2675.385, 9274.457),( 2690.403, 9300.469),( 2675.385, 9326.479),( 2675.385, 9673.518),( 2690.403, 9699.528),( 2675.385, 9725.539)), -- tube  84
    85 => (( 2705.420, 9274.457),( 2720.438, 9300.469),( 2705.420, 9326.479),( 2705.420, 9673.518),( 2720.438, 9699.528),( 2705.420, 9725.539)), -- tube  85
    86 => (( 2735.455, 9274.457),( 2750.472, 9300.469),( 2735.455, 9326.479),( 2735.455, 9673.518),( 2750.472, 9699.528),( 2735.455, 9725.539)), -- tube  86
    87 => (( 2765.490, 9274.457),( 2780.508, 9300.469),( 2765.490, 9326.479),( 2765.490, 9673.518),( 2780.508, 9699.528),( 2765.490, 9725.539)), -- tube  87
    88 => (( 2795.525, 9274.457),( 2810.542, 9300.469),( 2795.525, 9326.479),( 2795.525, 9673.518),( 2810.542, 9699.528),( 2795.525, 9725.539)), -- tube  88
    89 => (( 2825.560, 9274.457),( 2840.577, 9300.469),( 2825.560, 9326.479),( 2825.560, 9673.518),( 2840.577, 9699.528),( 2825.560, 9725.539)), -- tube  89
    90 => (( 2855.595, 9274.457),( 2870.613, 9300.469),( 2855.595, 9326.479),( 2855.595, 9673.518),( 2870.613, 9699.528),( 2855.595, 9725.539)), -- tube  90
    91 => (( 2885.630, 9274.457),( 2900.647, 9300.469),( 2885.630, 9326.479),( 2885.630, 9673.518),( 2900.647, 9699.528),( 2885.630, 9725.539)), -- tube  91
    92 => (( 2915.665, 9274.457),( 2930.683, 9300.469),( 2915.665, 9326.479),( 2915.665, 9673.518),( 2930.683, 9699.528),( 2915.665, 9725.539)), -- tube  92
    93 => (( 2945.700, 9274.457),( 2960.718, 9300.469),( 2945.700, 9326.479),( 2945.700, 9673.518),( 2960.718, 9699.528),( 2945.700, 9725.539)), -- tube  93
    94 => (( 2975.735, 9274.457),( 2990.752, 9300.469),( 2975.735, 9326.479),( 2975.735, 9673.518),( 2990.752, 9699.528),( 2975.735, 9725.539)), -- tube  94
    95 => (( 3005.735, 9274.457),( 3020.788, 9300.469),( 3005.770, 9326.479),( 3005.770, 9673.518),( 3020.788, 9699.528),( 3005.770, 9725.539)), -- tube  95
    96 => (( 3035.840, 9274.457),( 3050.857, 9300.469),( 3035.805, 9326.479),( 3035.805, 9673.518),( 3050.823, 9699.528),( 3035.805, 9725.539)), -- tube  96
    97 => (( 3065.840, 9274.457),( 3080.857, 9300.469),( 3065.840, 9326.479),( 3065.840, 9673.518),( 3080.857, 9699.528),( 3065.840, 9725.539)), -- tube  97
    98 => (( 3095.875, 9274.457),( 3110.893, 9300.469),( 3095.875, 9326.479),( 3095.875, 9673.518),( 3110.893, 9699.528),( 3095.875, 9725.539)), -- tube  98
    99 => (( 3125.910, 9274.457),( 3140.927, 9300.469),( 3125.910, 9326.479),( 3125.910, 9673.518),( 3140.927, 9699.528),( 3125.945, 9725.539)), -- tube  99
   100 => (( 3155.945, 9274.457),( 3170.962, 9300.469),( 3155.945, 9326.479),( 3155.945, 9673.518),( 3170.962, 9699.528),( 3155.945, 9725.539)), -- tube 100
   101 => (( 3185.980, 9274.457),( 3200.998, 9300.469),( 3185.980, 9326.479),( 3185.980, 9673.518),( 3200.998, 9699.528),( 3185.980, 9725.539)), -- tube 101
   102 => (( 3216.015, 9274.457),( 3231.032, 9300.469),( 3216.015, 9326.479),( 3216.015, 9673.518),( 3231.032, 9699.528),( 3216.015, 9725.539)), -- tube 102
   103 => (( 3246.050, 9274.457),( 3261.067, 9300.469),( 3246.050, 9326.479),( 3246.050, 9673.518),( 3261.067, 9699.528),( 3246.050, 9725.539)), -- tube 103
   104 => (( 3276.085, 9274.457),( 3291.103, 9300.469),( 3276.085, 9326.479),( 3276.085, 9673.518),( 3291.103, 9699.528),( 3276.085, 9725.539)), -- tube 104
   105 => (( 3306.120, 9274.457),( 3321.137, 9300.469),( 3306.120, 9326.479),( 3306.120, 9673.518),( 3321.137, 9699.528),( 3306.120, 9725.539)), -- tube 105
   106 => (( 3336.155, 9274.457),( 3351.173, 9300.469),( 3336.155, 9326.479),( 3336.155, 9673.518),( 3351.173, 9699.528),( 3336.155, 9725.539)), -- tube 106
   107 => (( 3366.190, 9274.457),( 3381.208, 9300.469),( 3366.190, 9326.479),( 3366.190, 9673.518),( 3381.208, 9699.528),( 3366.190, 9725.539)), -- tube 107
   108 => (( 3396.225, 9274.457),( 3411.242, 9300.469),( 3396.225, 9326.479),( 3396.225, 9673.518),( 3411.242, 9699.528),( 3396.225, 9725.539)), -- tube 108
   109 => (( 3426.260, 9274.457),( 3441.278, 9300.469),( 3426.260, 9326.479),( 3426.260, 9673.518),( 3441.278, 9699.528),( 3426.260, 9725.539)), -- tube 109
   110 => (( 3456.295, 9274.457),( 3471.312, 9300.469),( 3456.295, 9326.479),( 3456.295, 9673.518),( 3471.312, 9699.528),( 3456.295, 9725.539)), -- tube 110
   111 => (( 3486.330, 9274.457),( 3501.347, 9300.469),( 3486.330, 9326.479),( 3486.330, 9673.518),( 3501.383, 9699.528),( 3486.330, 9725.539)), -- tube 111
   112 => (( 3516.365, 9274.457),( 3531.383, 9300.469),( 3516.365, 9326.479),( 3516.365, 9673.518),( 3531.383, 9699.528),( 3516.365, 9725.539)), -- tube 112
   113 => (( 3546.400, 9274.457),( 3561.417, 9300.469),( 3546.400, 9326.479),( 3546.400, 9673.518),( 3561.417, 9699.528),( 3546.400, 9725.539)), -- tube 113
   114 => (( 3576.435, 9274.457),( 3591.452, 9300.469),( 3576.435, 9326.479),( 3576.435, 9673.518),( 3591.452, 9699.528),( 3576.435, 9725.539)), -- tube 114
   115 => (( 3606.470, 9274.457),( 3621.488, 9300.469),( 3606.470, 9326.479),( 3606.470, 9673.518),( 3621.488, 9699.528),( 3606.470, 9725.539)), -- tube 115
   116 => (( 3636.505, 9274.457),( 3651.522, 9300.469),( 3636.505, 9326.479),( 3636.505, 9673.518),( 3651.522, 9699.528),( 3636.505, 9725.539)), -- tube 116
   117 => (( 3666.540, 9274.457),( 3681.557, 9300.469),( 3666.540, 9326.479),( 3666.540, 9673.518),( 3681.557, 9699.528),( 3666.540, 9725.539)), -- tube 117
   118 => (( 3696.575, 9274.457),( 3711.593, 9300.469),( 3696.575, 9326.479),( 3696.575, 9673.518),( 3711.593, 9699.528),( 3696.575, 9725.539)), -- tube 118
   119 => (( 3726.610, 9274.457),( 3741.627, 9300.469),( 3726.610, 9326.479),( 3726.610, 9673.518),( 3741.627, 9699.528),( 3726.610, 9725.539)), -- tube 119
   120 => (( 3756.645, 9274.457),( 3771.663, 9300.469),( 3756.645, 9326.479),( 3756.645, 9673.518),( 3771.663, 9699.528),( 3756.645, 9725.539)), -- tube 120
   121 => (( 3786.680, 9274.457),( 3801.698, 9300.469),( 3786.680, 9326.479),( 3786.680, 9673.518),( 3801.698, 9699.528),( 3786.680, 9725.539)), -- tube 121
   122 => (( 3816.715, 9274.457),( 3831.732, 9300.469),( 3816.715, 9326.479),( 3816.715, 9673.518),( 3831.732, 9699.528),( 3816.715, 9725.539)), -- tube 122
   123 => (( 3846.750, 9274.457),( 3861.768, 9300.469),( 3846.750, 9326.479),( 3846.750, 9673.518),( 3861.768, 9699.528),( 3846.750, 9725.539)), -- tube 123
   124 => (( 3876.785, 9274.457),( 3891.802, 9300.469),( 3876.785, 9326.479),( 3876.785, 9673.518),( 3891.802, 9699.528),( 3876.785, 9725.539)), -- tube 124
   125 => (( 3906.820, 9274.457),( 3921.837, 9300.469),( 3906.820, 9326.479),( 3906.820, 9673.518),( 3921.837, 9699.528),( 3906.820, 9725.539)), -- tube 125
   126 => (( 3936.855, 9274.457),( 3951.873, 9300.469),( 3936.855, 9326.479),( 3936.855, 9673.518),( 3951.873, 9699.528),( 3936.855, 9725.539)), -- tube 126
   127 => (( 3966.890, 9274.457),( 3981.907, 9300.469),( 3966.890, 9326.479),( 3966.890, 9673.518),( 3981.907, 9699.528),( 3966.890, 9725.539)), -- tube 127
   128 => (( 3996.925, 9274.457),( 4011.942, 9300.469),( 3996.925, 9326.479),( 3996.925, 9673.518),( 4011.942, 9699.528),( 3996.925, 9725.539)), -- tube 128
   129 => (( 4026.960, 9274.457),( 4041.978, 9300.469),( 4026.960, 9326.479),( 4026.960, 9673.518),( 4041.978, 9699.528),( 4026.960, 9725.539)), -- tube 129
   130 => (( 4056.995, 9274.457),( 4072.012, 9300.469),( 4056.995, 9326.479),( 4056.995, 9673.518),( 4072.012, 9699.528),( 4056.995, 9725.539)), -- tube 130
   131 => (( 4087.030, 9274.457),( 4102.047, 9300.469),( 4087.030, 9326.479),( 4087.030, 9673.518),( 4102.047, 9699.528),( 4087.030, 9725.539)), -- tube 131
   132 => (( 4117.065, 9274.457),( 4132.083, 9300.469),( 4117.065, 9326.479),( 4117.065, 9673.518),( 4132.083, 9699.528),( 4117.065, 9725.539)), -- tube 132
   133 => (( 4147.100, 9274.457),( 4162.118, 9300.469),( 4147.100, 9326.479),( 4147.100, 9673.518),( 4162.118, 9699.528),( 4147.100, 9725.539)), -- tube 133
   134 => (( 4177.135, 9274.457),( 4192.152, 9300.469),( 4177.135, 9326.479),( 4177.135, 9673.518),( 4192.152, 9699.528),( 4177.135, 9725.539)), -- tube 134
   135 => (( 4207.170, 9274.457),( 4222.188, 9300.469),( 4207.170, 9326.479),( 4207.170, 9673.518),( 4222.188, 9699.528),( 4207.170, 9725.539)), -- tube 135
   136 => (( 4237.205, 9274.457),( 4252.223, 9300.469),( 4237.205, 9326.479),( 4237.205, 9673.518),( 4252.223, 9699.528),( 4237.205, 9725.539)), -- tube 136
   137 => (( 4267.240, 9274.457),( 4282.257, 9300.469),( 4267.240, 9326.479),( 4267.240, 9673.518),( 4282.257, 9699.528),( 4267.240, 9725.539)), -- tube 137
   138 => (( 4297.275, 9274.457),( 4312.292, 9300.469),( 4297.275, 9326.479),( 4297.275, 9673.518),( 4312.292, 9699.528),( 4297.275, 9725.539)), -- tube 138
   139 => (( 4327.310, 9274.457),( 4342.328, 9300.469),( 4327.310, 9326.479),( 4327.310, 9673.518),( 4342.328, 9699.528),( 4327.310, 9725.539)), -- tube 139
   140 => (( 4357.345, 9274.457),( 4372.362, 9300.469),( 4357.345, 9326.479),( 4357.345, 9673.518),( 4372.362, 9699.528),( 4357.345, 9725.539)), -- tube 140
   141 => (( 4387.380, 9274.457),( 4402.397, 9300.469),( 4387.380, 9326.479),( 4387.380, 9673.518),( 4402.397, 9699.528),( 4387.380, 9725.539)), -- tube 141
   142 => (( 4417.415, 9274.457),( 4432.433, 9300.469),( 4417.415, 9326.479),( 4417.415, 9673.518),( 4432.433, 9699.528),( 4417.415, 9725.539)), -- tube 142
   143 => (( 4447.450, 9274.457),( 4462.467, 9300.469),( 4447.450, 9326.479),( 4447.450, 9673.518),( 4462.467, 9699.528),( 4447.450, 9725.539)), -- tube 143
   144 => (( 4477.485, 9274.457),( 4492.502, 9300.469),( 4477.485, 9326.479),( 4477.485, 9673.518),( 4492.502, 9699.528),( 4477.485, 9725.539)), -- tube 144
   145 => (( 4525.000, 9274.457),( 4540.018, 9300.469),( 4525.000, 9326.479),( 4525.000, 9673.518),( 4540.018, 9699.528),( 4525.000, 9725.539)), -- tube 145
   146 => (( 4555.035, 9274.457),( 4570.053, 9300.469),( 4555.035, 9326.479),( 4555.035, 9673.518),( 4570.053, 9699.528),( 4555.035, 9725.539)), -- tube 146
   147 => (( 4585.070, 9274.457),( 4600.087, 9300.469),( 4585.070, 9326.479),( 4585.070, 9673.518),( 4600.087, 9699.528),( 4585.070, 9725.539)), -- tube 147
   148 => (( 4615.105, 9274.457),( 4630.123, 9300.469),( 4615.105, 9326.479),( 4615.105, 9673.518),( 4630.123, 9699.528),( 4615.105, 9725.539)), -- tube 148
   149 => (( 4645.140, 9274.457),( 4660.158, 9300.469),( 4645.140, 9326.479),( 4645.140, 9673.518),( 4660.158, 9699.528),( 4645.140, 9725.539)), -- tube 149
   150 => (( 4675.175, 9274.457),( 4690.192, 9300.469),( 4675.175, 9326.479),( 4675.175, 9673.518),( 4690.192, 9699.528),( 4675.175, 9725.539)), -- tube 150
   151 => (( 4705.210, 9274.457),( 4720.228, 9300.469),( 4705.210, 9326.479),( 4705.210, 9673.518),( 4720.228, 9699.528),( 4705.210, 9725.539)), -- tube 151
   152 => (( 4735.245, 9274.457),( 4750.263, 9300.469),( 4735.245, 9326.479),( 4735.245, 9673.518),( 4750.263, 9699.528),( 4735.245, 9725.539)), -- tube 152
   153 => (( 4765.280, 9274.457),( 4780.297, 9300.469),( 4765.280, 9326.479),( 4765.280, 9673.518),( 4780.297, 9699.528),( 4765.280, 9725.539)), -- tube 153
   154 => (( 4795.315, 9274.457),( 4810.333, 9300.469),( 4795.315, 9326.479),( 4795.315, 9673.518),( 4810.333, 9699.528),( 4795.315, 9725.539)), -- tube 154
   155 => (( 4825.350, 9274.457),( 4840.368, 9300.469),( 4825.350, 9326.479),( 4825.350, 9673.518),( 4840.368, 9699.528),( 4825.350, 9725.539)), -- tube 155
   156 => (( 4855.385, 9274.457),( 4870.402, 9300.469),( 4855.385, 9326.479),( 4855.385, 9673.518),( 4870.402, 9699.528),( 4855.385, 9725.539)), -- tube 156
   157 => (( 4885.420, 9274.457),( 4900.438, 9300.469),( 4885.420, 9326.479),( 4885.420, 9673.518),( 4900.438, 9699.528),( 4885.420, 9725.539)), -- tube 157
   158 => (( 4915.455, 9274.457),( 4930.473, 9300.469),( 4915.455, 9326.479),( 4915.455, 9673.518),( 4930.473, 9699.528),( 4915.455, 9725.539)), -- tube 158
   159 => (( 4945.490, 9274.457),( 4960.507, 9300.469),( 4945.490, 9326.479),( 4945.490, 9673.518),( 4960.507, 9699.528),( 4945.490, 9725.539)), -- tube 159
   160 => (( 4975.525, 9274.457),( 4990.542, 9300.469),( 4975.525, 9326.479),( 4975.525, 9673.518),( 4990.542, 9699.528),( 4975.525, 9725.539)), -- tube 160
   161 => (( 5005.560, 9274.457),( 5020.578, 9300.469),( 5005.560, 9326.479),( 5005.560, 9673.518),( 5020.578, 9699.528),( 5005.560, 9725.539)), -- tube 161
   162 => (( 5035.595, 9274.457),( 5050.612, 9300.469),( 5035.595, 9326.479),( 5035.595, 9673.518),( 5050.612, 9699.528),( 5035.595, 9725.539)), -- tube 162
   163 => (( 5065.630, 9274.457),( 5080.647, 9300.469),( 5065.630, 9326.479),( 5065.630, 9673.518),( 5080.647, 9699.528),( 5065.630, 9725.539)), -- tube 163
   164 => (( 5095.665, 9274.457),( 5110.683, 9300.469),( 5095.665, 9326.479),( 5095.665, 9673.518),( 5110.683, 9699.528),( 5095.665, 9725.539)), -- tube 164
   165 => (( 5125.700, 9274.457),( 5140.717, 9300.469),( 5125.700, 9326.479),( 5125.700, 9673.518),( 5140.717, 9699.528),( 5125.700, 9725.539)), -- tube 165
   166 => (( 5155.735, 9274.457),( 5170.752, 9300.469),( 5155.735, 9326.479),( 5155.735, 9673.518),( 5170.752, 9699.528),( 5155.735, 9725.539)), -- tube 166
   167 => (( 5185.770, 9274.457),( 5200.788, 9300.469),( 5185.770, 9326.479),( 5185.770, 9673.518),( 5200.788, 9699.528),( 5185.770, 9725.539)), -- tube 167
   168 => (( 5215.805, 9274.457),( 5230.822, 9300.469),( 5215.805, 9326.479),( 5215.805, 9673.518),( 5230.822, 9699.528),( 5215.805, 9725.539)), -- tube 168
   169 => (( 5245.840, 9274.457),( 5260.857, 9300.469),( 5245.840, 9326.479),( 5245.840, 9673.518),( 5260.857, 9699.528),( 5245.840, 9725.539)), -- tube 169
   170 => (( 5275.875, 9274.457),( 5290.893, 9300.469),( 5275.875, 9326.479),( 5275.875, 9673.518),( 5290.893, 9699.528),( 5275.875, 9725.539)), -- tube 170
   171 => (( 5305.910, 9274.457),( 5320.928, 9300.469),( 5305.910, 9326.479),( 5305.910, 9673.518),( 5320.928, 9699.528),( 5305.910, 9725.539)), -- tube 171
   172 => (( 5335.945, 9274.457),( 5350.962, 9300.469),( 5335.945, 9326.479),( 5335.945, 9673.518),( 5350.962, 9699.528),( 5335.945, 9725.539)), -- tube 172
   173 => (( 5365.980, 9274.457),( 5380.998, 9300.469),( 5365.980, 9326.479),( 5365.980, 9673.518),( 5380.998, 9699.528),( 5365.980, 9725.539)), -- tube 173
   174 => (( 5396.015, 9274.457),( 5411.033, 9300.469),( 5396.015, 9326.479),( 5396.015, 9673.518),( 5411.033, 9699.528),( 5396.015, 9725.539)), -- tube 174
   175 => (( 5426.050, 9274.457),( 5441.067, 9300.469),( 5426.050, 9326.479),( 5426.050, 9673.518),( 5441.067, 9699.528),( 5426.050, 9725.539)), -- tube 175
   176 => (( 5456.085, 9274.457),( 5471.103, 9300.469),( 5456.085, 9326.479),( 5456.085, 9673.518),( 5471.103, 9699.528),( 5456.085, 9725.539)), -- tube 176
   177 => (( 5486.120, 9274.457),( 5501.138, 9300.469),( 5486.120, 9326.479),( 5486.120, 9673.518),( 5501.138, 9699.528),( 5486.120, 9725.539)), -- tube 177
   178 => (( 5516.155, 9274.457),( 5531.172, 9300.469),( 5516.155, 9326.479),( 5516.155, 9673.518),( 5531.172, 9699.528),( 5516.155, 9725.539)), -- tube 178
   179 => (( 5546.190, 9274.457),( 5561.208, 9300.469),( 5546.190, 9326.479),( 5546.190, 9673.518),( 5561.208, 9699.528),( 5546.190, 9725.539)), -- tube 179
   180 => (( 5576.225, 9274.457),( 5591.243, 9300.469),( 5576.225, 9326.479),( 5576.225, 9673.518),( 5591.243, 9699.528),( 5576.225, 9725.539)), -- tube 180
   181 => (( 5606.260, 9274.457),( 5621.277, 9300.469),( 5606.260, 9326.479),( 5606.260, 9673.518),( 5621.277, 9699.528),( 5606.260, 9725.539)), -- tube 181
   182 => (( 5636.295, 9274.457),( 5651.312, 9300.469),( 5636.295, 9326.479),( 5636.295, 9673.518),( 5651.312, 9699.528),( 5636.295, 9725.539)), -- tube 182
   183 => (( 5666.330, 9274.457),( 5681.348, 9300.469),( 5666.330, 9326.479),( 5666.330, 9673.518),( 5681.348, 9699.528),( 5666.330, 9725.539)), -- tube 183
   184 => (( 5696.365, 9274.457),( 5711.382, 9300.469),( 5696.365, 9326.479),( 5696.365, 9673.518),( 5711.382, 9699.528),( 5696.365, 9725.539)), -- tube 184
   185 => (( 5726.400, 9274.457),( 5741.417, 9300.469),( 5726.400, 9326.479),( 5726.400, 9673.518),( 5741.417, 9699.528),( 5726.400, 9725.539)), -- tube 185
   186 => (( 5756.435, 9274.457),( 5771.453, 9300.469),( 5756.435, 9326.479),( 5756.435, 9673.518),( 5771.453, 9699.528),( 5756.435, 9725.539)), -- tube 186
   187 => (( 5786.470, 9274.457),( 5801.487, 9300.469),( 5786.470, 9326.479),( 5786.470, 9673.518),( 5801.487, 9699.528),( 5786.470, 9725.539)), -- tube 187
   188 => (( 5816.505, 9274.457),( 5831.522, 9300.469),( 5816.505, 9326.479),( 5816.505, 9673.518),( 5831.522, 9699.528),( 5816.505, 9725.539)), -- tube 188
   189 => (( 5846.540, 9274.457),( 5861.558, 9300.469),( 5846.540, 9326.479),( 5846.540, 9673.518),( 5861.558, 9699.528),( 5846.540, 9725.539)), -- tube 189
   190 => (( 5876.575, 9274.457),( 5891.592, 9300.469),( 5876.575, 9326.479),( 5876.575, 9673.518),( 5891.592, 9699.528),( 5876.575, 9725.539)), -- tube 190
   191 => (( 5906.610, 9274.457),( 5921.627, 9300.469),( 5906.610, 9326.479),( 5906.610, 9673.518),( 5921.627, 9699.528),( 5906.610, 9725.539)), -- tube 191
   192 => (( 5936.645, 9274.457),( 5951.663, 9300.469),( 5936.645, 9326.479),( 5936.645, 9673.518),( 5951.663, 9699.528),( 5936.645, 9725.539)), -- tube 192
   193 => (( 5966.680, 9274.457),( 5981.697, 9300.469),( 5966.680, 9326.479),( 5966.680, 9673.518),( 5981.697, 9699.528),( 5966.680, 9725.539)), -- tube 193
   194 => (( 5996.715, 9274.457),( 6011.732, 9300.469),( 5996.715, 9326.479),( 5996.715, 9673.518),( 6011.732, 9699.528),( 5996.715, 9725.539)), -- tube 194
   195 => (( 6026.750, 9274.457),( 6041.768, 9300.469),( 6026.750, 9326.479),( 6026.750, 9673.518),( 6041.768, 9699.528),( 6026.750, 9725.539)), -- tube 195
   196 => (( 6056.785, 9274.457),( 6071.803, 9300.469),( 6056.785, 9326.479),( 6056.785, 9673.518),( 6071.803, 9699.528),( 6056.785, 9725.539)), -- tube 196
   197 => (( 6086.820, 9274.457),( 6101.837, 9300.469),( 6086.820, 9326.479),( 6086.820, 9673.518),( 6101.837, 9699.528),( 6086.820, 9725.539)), -- tube 197
   198 => (( 6116.855, 9274.457),( 6131.873, 9300.469),( 6116.855, 9326.479),( 6116.855, 9673.518),( 6131.873, 9699.528),( 6116.855, 9725.539)), -- tube 198
   199 => (( 6146.890, 9274.457),( 6161.908, 9300.469),( 6146.890, 9326.479),( 6146.890, 9673.518),( 6161.908, 9699.528),( 6146.890, 9725.539)), -- tube 199
   200 => (( 6176.925, 9274.457),( 6191.942, 9300.469),( 6176.925, 9326.479),( 6176.925, 9673.518),( 6191.942, 9699.528),( 6176.925, 9725.539)), -- tube 200
   201 => (( 6225.000, 9274.457),( 6240.018, 9300.469),( 6225.000, 9326.479),( 6225.000, 9673.518),( 6240.018, 9699.528),( 6225.000, 9725.539)), -- tube 201
   202 => (( 6255.035, 9274.457),( 6270.053, 9300.469),( 6255.035, 9326.479),( 6255.035, 9673.518),( 6270.053, 9699.528),( 6255.035, 9725.539)), -- tube 202
   203 => (( 6285.070, 9274.457),( 6300.087, 9300.469),( 6285.070, 9326.479),( 6285.070, 9673.518),( 6300.087, 9699.528),( 6285.070, 9725.539)), -- tube 203
   204 => (( 6315.105, 9274.457),( 6330.123, 9300.469),( 6315.105, 9326.479),( 6315.105, 9673.518),( 6330.123, 9699.528),( 6315.105, 9725.539)), -- tube 204
   205 => (( 6345.140, 9274.457),( 6360.158, 9300.469),( 6345.140, 9326.479),( 6345.140, 9673.518),( 6360.158, 9699.528),( 6345.140, 9725.539)), -- tube 205
   206 => (( 6375.175, 9274.457),( 6390.192, 9300.469),( 6375.175, 9326.479),( 6375.175, 9673.518),( 6390.192, 9699.528),( 6375.175, 9725.539)), -- tube 206
   207 => (( 6405.210, 9274.457),( 6420.228, 9300.469),( 6405.210, 9326.479),( 6405.210, 9673.518),( 6420.228, 9699.528),( 6405.210, 9725.539)), -- tube 207
   208 => (( 6435.245, 9274.457),( 6450.263, 9300.469),( 6435.245, 9326.479),( 6435.245, 9673.518),( 6450.263, 9699.528),( 6435.245, 9725.539)), -- tube 208
   209 => (( 6465.280, 9274.457),( 6480.297, 9300.469),( 6465.280, 9326.479),( 6465.280, 9673.518),( 6480.297, 9699.528),( 6465.280, 9725.539)), -- tube 209
   210 => (( 6495.315, 9274.457),( 6510.333, 9300.469),( 6495.315, 9326.479),( 6495.315, 9673.518),( 6510.333, 9699.528),( 6495.315, 9725.539)), -- tube 210
   211 => (( 6525.350, 9274.457),( 6540.368, 9300.469),( 6525.350, 9326.479),( 6525.350, 9673.518),( 6540.368, 9699.528),( 6525.350, 9725.539)), -- tube 211
   212 => (( 6555.385, 9274.457),( 6570.402, 9300.469),( 6555.385, 9326.479),( 6555.385, 9673.518),( 6570.402, 9699.528),( 6555.385, 9725.539)), -- tube 212
   213 => (( 6585.420, 9274.457),( 6600.438, 9300.469),( 6585.420, 9326.479),( 6585.420, 9673.518),( 6600.438, 9699.528),( 6585.420, 9725.539)), -- tube 213
   214 => (( 6615.455, 9274.457),( 6630.473, 9300.469),( 6615.455, 9326.479),( 6615.455, 9673.518),( 6630.473, 9699.528),( 6615.455, 9725.539)), -- tube 214
   215 => (( 6645.490, 9274.457),( 6660.507, 9300.469),( 6645.490, 9326.479),( 6645.490, 9673.518),( 6660.507, 9699.528),( 6645.490, 9725.539)), -- tube 215
   216 => (( 6675.525, 9274.457),( 6690.542, 9300.469),( 6675.525, 9326.479),( 6675.525, 9673.518),( 6690.542, 9699.528),( 6675.525, 9725.539)), -- tube 216
   217 => (( 6705.560, 9274.457),( 6720.578, 9300.469),( 6705.560, 9326.479),( 6705.560, 9673.518),( 6720.578, 9699.528),( 6705.560, 9725.539)), -- tube 217
   218 => (( 6735.595, 9274.457),( 6750.612, 9300.469),( 6735.595, 9326.479),( 6735.595, 9673.518),( 6750.612, 9699.528),( 6735.595, 9725.539)), -- tube 218
   219 => (( 6765.630, 9274.457),( 6780.647, 9300.469),( 6765.630, 9326.479),( 6765.630, 9673.518),( 6780.647, 9699.528),( 6765.630, 9725.539)), -- tube 219
   220 => (( 6795.665, 9274.457),( 6810.683, 9300.469),( 6795.665, 9326.479),( 6795.665, 9673.518),( 6810.683, 9699.528),( 6795.665, 9725.539)), -- tube 220
   221 => (( 6825.700, 9274.457),( 6840.717, 9300.469),( 6825.700, 9326.479),( 6825.700, 9673.518),( 6840.717, 9699.528),( 6825.700, 9725.539)), -- tube 221
   222 => (( 6855.735, 9274.457),( 6870.752, 9300.469),( 6855.735, 9326.479),( 6855.735, 9673.518),( 6870.752, 9699.528),( 6855.735, 9725.539)), -- tube 222
   223 => (( 6885.770, 9274.457),( 6900.788, 9300.469),( 6885.770, 9326.479),( 6885.770, 9673.518),( 6900.788, 9699.528),( 6885.770, 9725.539)), -- tube 223
   224 => (( 6915.805, 9274.457),( 6930.822, 9300.469),( 6915.805, 9326.479),( 6915.805, 9673.518),( 6930.822, 9699.528),( 6915.805, 9725.539)), -- tube 224
   225 => (( 6945.840, 9274.457),( 6960.857, 9300.469),( 6945.840, 9326.479),( 6945.840, 9673.518),( 6960.857, 9699.528),( 6945.840, 9725.539)), -- tube 225
   226 => (( 6975.875, 9274.457),( 6990.893, 9300.469),( 6975.875, 9326.479),( 6975.875, 9673.518),( 6990.893, 9699.528),( 6975.875, 9725.539)), -- tube 226
   227 => (( 7005.910, 9274.457),( 7020.928, 9300.469),( 7005.910, 9326.479),( 7005.910, 9673.518),( 7020.928, 9699.528),( 7005.910, 9725.539)), -- tube 227
   228 => (( 7035.945, 9274.457),( 7050.962, 9300.469),( 7035.945, 9326.479),( 7035.945, 9673.518),( 7050.962, 9699.528),( 7035.945, 9725.539)), -- tube 228
   229 => (( 7065.980, 9274.457),( 7080.998, 9300.469),( 7065.980, 9326.479),( 7065.980, 9673.518),( 7080.998, 9699.528),( 7065.980, 9725.539)), -- tube 229
   230 => (( 7096.015, 9274.457),( 7111.033, 9300.469),( 7096.015, 9326.479),( 7096.015, 9673.518),( 7111.033, 9699.528),( 7096.015, 9725.539)), -- tube 230
   231 => (( 7126.050, 9274.457),( 7141.067, 9300.469),( 7126.050, 9326.479),( 7126.050, 9673.518),( 7141.067, 9699.528),( 7126.050, 9725.539)), -- tube 231
   232 => (( 7156.085, 9274.457),( 7171.103, 9300.469),( 7156.085, 9326.479),( 7156.085, 9673.518),( 7171.103, 9699.528),( 7156.085, 9725.539)), -- tube 232
   233 => (( 7186.120, 9274.457),( 7201.138, 9300.469),( 7186.120, 9326.479),( 7186.120, 9673.518),( 7201.138, 9699.528),( 7186.120, 9725.539)), -- tube 233
   234 => (( 7216.155, 9274.457),( 7231.172, 9300.469),( 7216.155, 9326.479),( 7216.155, 9673.518),( 7231.172, 9699.528),( 7216.155, 9725.539)), -- tube 234
   235 => (( 7246.190, 9274.457),( 7261.208, 9300.469),( 7246.190, 9326.479),( 7246.190, 9673.518),( 7261.208, 9699.528),( 7246.190, 9725.539)), -- tube 235
   236 => (( 7276.225, 9274.457),( 7291.243, 9300.469),( 7276.225, 9326.479),( 7276.225, 9673.518),( 7291.243, 9699.528),( 7276.225, 9725.539)), -- tube 236
   237 => (( 7306.260, 9274.457),( 7321.277, 9300.469),( 7306.260, 9326.479),( 7306.260, 9673.518),( 7321.277, 9699.528),( 7306.260, 9725.539)), -- tube 237
   238 => (( 7336.295, 9274.457),( 7351.312, 9300.469),( 7336.295, 9326.479),( 7336.295, 9673.518),( 7351.312, 9699.528),( 7336.295, 9725.539)), -- tube 238
   239 => (( 7366.330, 9274.457),( 7381.348, 9300.469),( 7366.330, 9326.479),( 7366.330, 9673.518),( 7381.348, 9699.528),( 7366.330, 9725.539)), -- tube 239
   240 => (( 7396.365, 9274.457),( 7411.382, 9300.469),( 7396.365, 9326.479),( 7396.365, 9673.518),( 7411.382, 9699.528),( 7396.365, 9725.539)), -- tube 240
   241 => (( 7426.400, 9274.457),( 7441.417, 9300.469),( 7426.400, 9326.479),( 7426.400, 9673.518),( 7441.417, 9699.528),( 7426.400, 9725.539)), -- tube 241
   242 => (( 7456.435, 9274.457),( 7471.453, 9300.469),( 7456.435, 9326.479),( 7456.435, 9673.518),( 7471.453, 9699.528),( 7456.435, 9725.539)), -- tube 242
   243 => (( 7486.470, 9274.457),( 7501.487, 9300.469),( 7486.470, 9326.479),( 7486.470, 9673.518),( 7501.487, 9699.528),( 7486.470, 9725.539)), -- tube 243
   244 => (( 7516.505, 9274.457),( 7531.522, 9300.469),( 7516.505, 9326.479),( 7516.505, 9673.518),( 7531.522, 9699.528),( 7516.505, 9725.539)), -- tube 244
   245 => (( 7546.540, 9274.457),( 7561.558, 9300.469),( 7546.540, 9326.479),( 7546.540, 9673.518),( 7561.558, 9699.528),( 7546.540, 9725.539)), -- tube 245
   246 => (( 7576.575, 9274.457),( 7591.592, 9300.469),( 7576.575, 9326.479),( 7576.575, 9673.518),( 7591.592, 9699.528),( 7576.575, 9725.539)), -- tube 246
   247 => (( 7606.610, 9274.457),( 7621.627, 9300.469),( 7606.610, 9326.479),( 7606.610, 9673.518),( 7621.627, 9699.528),( 7606.610, 9725.539)), -- tube 247
   248 => (( 7636.645, 9274.457),( 7651.663, 9300.469),( 7636.645, 9326.479),( 7636.645, 9673.518),( 7651.663, 9699.528),( 7636.645, 9725.539)), -- tube 248
   249 => (( 7666.680, 9274.457),( 7681.697, 9300.469),( 7666.680, 9326.479),( 7666.680, 9673.518),( 7681.697, 9699.528),( 7666.680, 9725.539)), -- tube 249
   250 => (( 7696.715, 9274.457),( 7711.732, 9300.469),( 7696.715, 9326.479),( 7696.715, 9673.518),( 7711.732, 9699.528),( 7696.715, 9725.539)), -- tube 250
   251 => (( 7726.750, 9274.457),( 7741.768, 9300.469),( 7726.750, 9326.479),( 7726.750, 9673.518),( 7741.768, 9699.528),( 7726.750, 9725.539)), -- tube 251
   252 => (( 7756.785, 9274.457),( 7771.803, 9300.469),( 7756.785, 9326.479),( 7756.785, 9673.518),( 7771.803, 9699.528),( 7756.785, 9725.539)), -- tube 252
   253 => (( 7786.820, 9274.457),( 7801.837, 9300.469),( 7786.820, 9326.479),( 7786.820, 9673.518),( 7801.837, 9699.528),( 7786.820, 9725.539)), -- tube 253
   254 => (( 7816.855, 9274.457),( 7831.873, 9300.469),( 7816.855, 9326.479),( 7816.855, 9673.518),( 7831.873, 9699.528),( 7816.855, 9725.539)), -- tube 254
   255 => (( 7846.890, 9274.457),( 7861.908, 9300.469),( 7846.890, 9326.479),( 7846.890, 9673.518),( 7861.908, 9699.528),( 7846.890, 9725.539)), -- tube 255
   256 => (( 7876.925, 9274.457),( 7891.942, 9300.469),( 7876.925, 9326.479),( 7876.925, 9673.518),( 7891.942, 9699.528),( 7876.925, 9725.539)), -- tube 256
   257 => (( 7906.960, 9274.457),( 7921.978, 9300.469),( 7906.960, 9326.479),( 7906.960, 9673.518),( 7921.978, 9699.528),( 7906.960, 9725.539)), -- tube 257
   258 => (( 7936.995, 9274.457),( 7952.013, 9300.469),( 7936.995, 9326.479),( 7936.995, 9673.518),( 7952.013, 9699.528),( 7936.995, 9725.539)), -- tube 258
   259 => (( 7967.030, 9274.457),( 7982.047, 9300.469),( 7967.030, 9326.479),( 7967.030, 9673.518),( 7982.047, 9699.528),( 7967.030, 9725.539)), -- tube 259
   260 => (( 7997.065, 9274.457),( 8012.083, 9300.469),( 7997.065, 9326.479),( 7997.065, 9673.518),( 8012.083, 9699.528),( 7997.065, 9725.539)), -- tube 260
   261 => (( 8027.100, 9274.457),( 8042.118, 9300.469),( 8027.100, 9326.479),( 8027.100, 9673.518),( 8042.118, 9699.528),( 8027.100, 9725.539)), -- tube 261
   262 => (( 8057.135, 9274.457),( 8072.152, 9300.469),( 8057.135, 9326.479),( 8057.135, 9673.518),( 8072.152, 9699.528),( 8057.135, 9725.539)), -- tube 262
   263 => (( 8087.170, 9274.457),( 8102.188, 9300.469),( 8087.170, 9326.479),( 8087.170, 9673.518),( 8102.188, 9699.528),( 8087.170, 9725.539)), -- tube 263
   264 => (( 8117.205, 9274.457),( 8132.223, 9300.469),( 8117.205, 9326.479),( 8117.205, 9673.518),( 8132.223, 9699.528),( 8117.205, 9725.539)), -- tube 264
   265 => (( 8147.240, 9274.457),( 8162.257, 9300.469),( 8147.240, 9326.479),( 8147.240, 9673.518),( 8162.257, 9699.528),( 8147.240, 9725.539)), -- tube 265
   266 => (( 8177.275, 9274.457),( 8192.293, 9300.469),( 8177.275, 9326.479),( 8177.275, 9673.518),( 8192.293, 9699.528),( 8177.275, 9725.539)), -- tube 266
   267 => (( 8207.310, 9274.457),( 8222.327, 9300.469),( 8207.310, 9326.479),( 8207.310, 9673.518),( 8222.327, 9699.528),( 8207.310, 9725.539)), -- tube 267
   268 => (( 8237.345, 9274.457),( 8252.362, 9300.469),( 8237.345, 9326.479),( 8237.345, 9673.518),( 8252.362, 9699.528),( 8237.345, 9725.539)), -- tube 268
   269 => (( 8267.380, 9274.457),( 8282.397, 9300.469),( 8267.380, 9326.479),( 8267.380, 9673.518),( 8282.397, 9699.528),( 8267.380, 9725.539)), -- tube 269
   270 => (( 8297.415, 9274.457),( 8312.433, 9300.469),( 8297.415, 9326.479),( 8297.415, 9673.518),( 8312.433, 9699.528),( 8297.415, 9725.539)), -- tube 270
   271 => (( 8327.450, 9274.457),( 8342.468, 9300.469),( 8327.450, 9326.479),( 8327.450, 9673.518),( 8342.468, 9699.528),( 8327.450, 9725.539)), -- tube 271
   272 => (( 8357.485, 9274.457),( 8372.503, 9300.469),( 8357.485, 9326.479),( 8357.485, 9673.518),( 8372.503, 9699.528),( 8357.485, 9725.539)), -- tube 272
   273 => (( 8405.000, 9274.457),( 8420.018, 9300.469),( 8405.000, 9326.479),( 8405.000, 9673.518),( 8420.018, 9699.528),( 8405.000, 9725.539)), -- tube 273
   274 => (( 8435.035, 9274.457),( 8450.053, 9300.469),( 8435.035, 9326.479),( 8435.035, 9673.518),( 8450.053, 9699.528),( 8435.035, 9725.539)), -- tube 274
   275 => (( 8465.070, 9274.457),( 8480.088, 9300.469),( 8465.070, 9326.479),( 8465.070, 9673.518),( 8480.088, 9699.528),( 8465.070, 9725.539)), -- tube 275
   276 => (( 8495.105, 9274.457),( 8510.122, 9300.469),( 8495.105, 9326.479),( 8495.105, 9673.518),( 8510.122, 9699.528),( 8495.105, 9725.539)), -- tube 276
   277 => (( 8525.140, 9274.457),( 8540.157, 9300.469),( 8525.140, 9326.479),( 8525.140, 9673.518),( 8540.157, 9699.528),( 8525.140, 9725.539)), -- tube 277
   278 => (( 8555.175, 9274.457),( 8570.192, 9300.469),( 8555.175, 9326.479),( 8555.175, 9673.518),( 8570.192, 9699.528),( 8555.175, 9725.539)), -- tube 278
   279 => (( 8585.210, 9274.457),( 8600.228, 9300.469),( 8585.210, 9326.479),( 8585.210, 9673.518),( 8600.228, 9699.528),( 8585.210, 9725.539)), -- tube 279
   280 => (( 8615.245, 9274.457),( 8630.263, 9300.469),( 8615.245, 9326.479),( 8615.245, 9673.518),( 8630.263, 9699.528),( 8615.245, 9725.539)), -- tube 280
   281 => (( 8645.280, 9274.457),( 8660.298, 9300.469),( 8645.280, 9326.479),( 8645.280, 9673.518),( 8660.298, 9699.528),( 8645.280, 9725.539)), -- tube 281
   282 => (( 8675.315, 9274.457),( 8690.332, 9300.469),( 8675.315, 9326.479),( 8675.315, 9673.518),( 8690.332, 9699.528),( 8675.315, 9725.539)), -- tube 282
   283 => (( 8705.350, 9274.457),( 8720.367, 9300.469),( 8705.350, 9326.479),( 8705.350, 9673.518),( 8720.367, 9699.528),( 8705.350, 9725.539)), -- tube 283
   284 => (( 8735.385, 9274.457),( 8750.402, 9300.469),( 8735.385, 9326.479),( 8735.385, 9673.518),( 8750.402, 9699.528),( 8735.385, 9725.539)), -- tube 284
   285 => (( 8765.420, 9274.457),( 8780.438, 9300.469),( 8765.420, 9326.479),( 8765.420, 9673.518),( 8780.438, 9699.528),( 8765.420, 9725.539)), -- tube 285
   286 => (( 8795.455, 9274.457),( 8810.473, 9300.469),( 8795.455, 9326.479),( 8795.455, 9673.518),( 8810.473, 9699.528),( 8795.455, 9725.539)), -- tube 286
   287 => (( 8825.490, 9274.457),( 8840.508, 9300.469),( 8825.490, 9326.479),( 8825.490, 9673.518),( 8840.508, 9699.528),( 8825.490, 9725.539)), -- tube 287
   288 => (( 8855.525, 9274.457),( 8870.543, 9300.469),( 8855.525, 9326.479),( 8855.525, 9673.518),( 8870.543, 9699.528),( 8855.525, 9725.539)), -- tube 288
   289 => (( 8885.560, 9274.457),( 8900.577, 9300.469),( 8885.560, 9326.479),( 8885.560, 9673.518),( 8900.577, 9699.528),( 8885.560, 9725.539)), -- tube 289
   290 => (( 8915.595, 9274.457),( 8930.612, 9300.469),( 8915.595, 9326.479),( 8915.595, 9673.518),( 8930.612, 9699.528),( 8915.595, 9725.539)), -- tube 290
   291 => (( 8945.630, 9274.457),( 8960.647, 9300.469),( 8945.630, 9326.479),( 8945.630, 9673.518),( 8960.647, 9699.528),( 8945.630, 9725.539)), -- tube 291
   292 => (( 8975.665, 9274.457),( 8990.683, 9300.469),( 8975.665, 9326.479),( 8975.665, 9673.518),( 8990.683, 9699.528),( 8975.665, 9725.539)), -- tube 292
   293 => (( 9005.700, 9274.457),( 9020.718, 9300.469),( 9005.700, 9326.479),( 9005.700, 9673.518),( 9020.718, 9699.528),( 9005.700, 9725.539)), -- tube 293
   294 => (( 9035.735, 9274.457),( 9050.753, 9300.469),( 9035.735, 9326.479),( 9035.735, 9673.518),( 9050.753, 9699.528),( 9035.735, 9725.539)), -- tube 294
   295 => (( 9065.770, 9274.457),( 9080.787, 9300.469),( 9065.770, 9326.479),( 9065.770, 9673.518),( 9080.787, 9699.528),( 9065.770, 9725.539)), -- tube 295
   296 => (( 9095.805, 9274.457),( 9110.822, 9300.469),( 9095.805, 9326.479),( 9095.805, 9673.518),( 9110.822, 9699.528),( 9095.805, 9725.539)), -- tube 296
   297 => (( 9125.840, 9274.457),( 9140.857, 9300.469),( 9125.840, 9326.479),( 9125.840, 9673.518),( 9140.857, 9699.528),( 9125.840, 9725.539)), -- tube 297
   298 => (( 9155.875, 9274.457),( 9170.893, 9300.469),( 9155.875, 9326.479),( 9155.875, 9673.518),( 9170.893, 9699.528),( 9155.875, 9725.539)), -- tube 298
   299 => (( 9185.910, 9274.457),( 9200.928, 9300.469),( 9185.910, 9326.479),( 9185.910, 9673.518),( 9200.928, 9699.528),( 9185.910, 9725.539)), -- tube 299
   300 => (( 9215.945, 9274.457),( 9230.963, 9300.469),( 9215.945, 9326.479),( 9215.945, 9673.518),( 9230.963, 9699.528),( 9215.945, 9725.539)), -- tube 300
   301 => (( 9245.980, 9274.457),( 9260.997, 9300.469),( 9245.980, 9326.479),( 9245.980, 9673.518),( 9260.997, 9699.528),( 9245.980, 9725.539)), -- tube 301
   302 => (( 9276.015, 9274.457),( 9291.032, 9300.469),( 9276.015, 9326.479),( 9276.015, 9673.518),( 9291.032, 9699.528),( 9276.015, 9725.539)), -- tube 302
   303 => (( 9306.050, 9274.457),( 9321.067, 9300.469),( 9306.050, 9326.479),( 9306.050, 9673.518),( 9321.067, 9699.528),( 9306.050, 9725.539)), -- tube 303
   304 => (( 9336.085, 9274.457),( 9351.103, 9300.469),( 9336.085, 9326.479),( 9336.085, 9673.518),( 9351.103, 9699.528),( 9336.085, 9725.539)), -- tube 304
   305 => (( 9366.120, 9274.457),( 9381.138, 9300.469),( 9366.120, 9326.479),( 9366.120, 9673.518),( 9381.138, 9699.528),( 9366.120, 9725.539)), -- tube 305
   306 => (( 9396.155, 9274.457),( 9411.173, 9300.469),( 9396.155, 9326.479),( 9396.155, 9673.518),( 9411.173, 9699.528),( 9396.155, 9725.539)), -- tube 306
   307 => (( 9426.190, 9274.457),( 9441.207, 9300.469),( 9426.190, 9326.479),( 9426.190, 9673.518),( 9441.207, 9699.528),( 9426.190, 9725.539)), -- tube 307
   308 => (( 9456.225, 9274.457),( 9471.242, 9300.469),( 9456.225, 9326.479),( 9456.225, 9673.518),( 9471.242, 9699.528),( 9456.225, 9725.539)), -- tube 308
   309 => (( 9486.260, 9274.457),( 9501.277, 9300.469),( 9486.260, 9326.479),( 9486.260, 9673.518),( 9501.277, 9699.528),( 9486.260, 9725.539)), -- tube 309
   310 => (( 9516.295, 9274.457),( 9531.312, 9300.469),( 9516.295, 9326.479),( 9516.295, 9673.518),( 9531.312, 9699.528),( 9516.295, 9725.539)), -- tube 310
   311 => (( 9546.330, 9274.457),( 9561.348, 9300.469),( 9546.330, 9326.479),( 9546.330, 9673.518),( 9561.348, 9699.528),( 9546.330, 9725.539)), -- tube 311
   312 => (( 9576.365, 9274.457),( 9591.383, 9300.469),( 9576.365, 9326.479),( 9576.365, 9673.518),( 9591.383, 9699.528),( 9576.365, 9725.539)), -- tube 312
   313 => (( 9606.400, 9274.457),( 9621.418, 9300.469),( 9606.400, 9326.479),( 9606.400, 9673.518),( 9621.418, 9699.528),( 9606.400, 9725.539)), -- tube 313
   314 => (( 9636.435, 9274.457),( 9651.452, 9300.469),( 9636.435, 9326.479),( 9636.435, 9673.518),( 9651.452, 9699.528),( 9636.435, 9725.539)), -- tube 314
   315 => (( 9666.470, 9274.457),( 9681.487, 9300.469),( 9666.470, 9326.479),( 9666.470, 9673.518),( 9681.487, 9699.528),( 9666.470, 9725.539)), -- tube 315
   316 => (( 9696.505, 9274.457),( 9711.522, 9300.469),( 9696.505, 9326.479),( 9696.505, 9673.518),( 9711.522, 9699.528),( 9696.505, 9725.539)), -- tube 316
   317 => (( 9726.540, 9274.457),( 9741.558, 9300.469),( 9726.540, 9326.479),( 9726.540, 9673.518),( 9741.558, 9699.528),( 9726.540, 9725.539)), -- tube 317
   318 => (( 9756.575, 9274.457),( 9771.593, 9300.469),( 9756.575, 9326.479),( 9756.575, 9673.518),( 9771.593, 9699.528),( 9756.575, 9725.539)), -- tube 318
   319 => (( 9786.610, 9274.457),( 9801.628, 9300.469),( 9786.610, 9326.479),( 9786.610, 9673.518),( 9801.628, 9699.528),( 9786.610, 9725.539)), -- tube 319
   320 => (( 9816.645, 9274.457),( 9831.662, 9300.469),( 9816.645, 9326.479),( 9816.645, 9673.518),( 9831.662, 9699.528),( 9816.645, 9725.539)), -- tube 320
   321 => (( 9846.680, 9274.457),( 9861.697, 9300.469),( 9846.680, 9326.479),( 9846.680, 9673.518),( 9861.697, 9699.528),( 9846.680, 9725.539)), -- tube 321
   322 => (( 9876.715, 9274.457),( 9891.732, 9300.469),( 9876.715, 9326.479),( 9876.715, 9673.518),( 9891.732, 9699.528),( 9876.715, 9725.539)), -- tube 322
   323 => (( 9906.750, 9274.457),( 9921.768, 9300.469),( 9906.750, 9326.479),( 9906.750, 9673.518),( 9921.768, 9699.528),( 9906.750, 9725.539)), -- tube 323
   324 => (( 9936.785, 9274.457),( 9951.803, 9300.469),( 9936.785, 9326.479),( 9936.785, 9673.518),( 9951.803, 9699.528),( 9936.785, 9725.539)), -- tube 324
   325 => (( 9966.820, 9274.457),( 9981.838, 9300.469),( 9966.820, 9326.479),( 9966.820, 9673.518),( 9981.838, 9699.528),( 9966.820, 9725.539)), -- tube 325
   326 => (( 9996.855, 9274.457),(10011.872, 9300.469),( 9996.855, 9326.479),( 9996.855, 9673.518),(10011.872, 9699.528),( 9996.855, 9725.539)), -- tube 326
   327 => ((10026.890, 9274.457),(10041.907, 9300.469),(10026.890, 9326.479),(10026.890, 9673.518),(10041.907, 9699.528),(10026.890, 9725.539)), -- tube 327
   328 => ((10056.925, 9274.457),(10071.942, 9300.469),(10056.925, 9326.479),(10056.925, 9673.518),(10071.942, 9699.528),(10056.925, 9725.539)), -- tube 328
   329 => ((10086.960, 9274.457),(10101.978, 9300.469),(10086.960, 9326.479),(10086.960, 9673.518),(10101.978, 9699.528),(10086.960, 9725.539)), -- tube 329
   330 => ((10116.995, 9274.457),(10132.013, 9300.469),(10116.995, 9326.479),(10116.995, 9673.518),(10132.013, 9699.528),(10116.995, 9725.539)), -- tube 330
   331 => ((10147.030, 9274.457),(10162.048, 9300.469),(10147.030, 9326.479),(10147.030, 9673.518),(10162.048, 9699.528),(10147.030, 9725.539)), -- tube 331
   332 => ((10177.065, 9274.457),(10192.082, 9300.469),(10177.065, 9326.479),(10177.065, 9673.518),(10192.082, 9699.528),(10177.065, 9725.539)), -- tube 332
   333 => ((10207.100, 9274.457),(10222.117, 9300.469),(10207.100, 9326.479),(10207.100, 9673.518),(10222.117, 9699.528),(10207.100, 9725.539)), -- tube 333
   334 => ((10237.135, 9274.457),(10252.152, 9300.469),(10237.135, 9326.479),(10237.135, 9673.518),(10252.152, 9699.528),(10237.135, 9725.539)), -- tube 334
   335 => ((10267.170, 9274.457),(10282.188, 9300.469),(10267.170, 9326.479),(10267.170, 9673.518),(10282.188, 9699.528),(10267.170, 9725.539)), -- tube 335
   336 => ((10297.205, 9274.457),(10312.223, 9300.469),(10297.205, 9326.479),(10297.205, 9673.518),(10312.223, 9699.528),(10297.205, 9725.539)), -- tube 336
   337 => ((10327.240, 9274.457),(10342.258, 9300.469),(10327.240, 9326.479),(10327.240, 9673.518),(10342.258, 9699.528),(10327.240, 9725.539)), -- tube 337
   338 => ((10357.275, 9274.457),(10372.293, 9300.469),(10357.275, 9326.479),(10357.275, 9673.518),(10372.293, 9699.528),(10357.275, 9725.539)), -- tube 338
   339 => ((10387.310, 9274.457),(10402.327, 9300.469),(10387.310, 9326.479),(10387.310, 9673.518),(10402.327, 9699.528),(10387.310, 9725.539)), -- tube 339
   340 => ((10417.345, 9274.457),(10432.362, 9300.469),(10417.345, 9326.479),(10417.345, 9673.518),(10432.362, 9699.528),(10417.345, 9725.539)), -- tube 340
   341 => ((10447.380, 9274.457),(10462.397, 9300.469),(10447.380, 9326.479),(10447.380, 9673.518),(10462.397, 9699.528),(10447.380, 9725.539)), -- tube 341
   342 => ((10477.415, 9274.457),(10492.433, 9300.469),(10477.415, 9326.479),(10477.415, 9673.518),(10492.433, 9699.528),(10477.415, 9725.539)), -- tube 342
   343 => ((10507.450, 9274.457),(10522.468, 9300.469),(10507.450, 9326.479),(10507.450, 9673.518),(10522.468, 9699.528),(10507.450, 9725.539)), -- tube 343
   344 => ((10537.485, 9274.457),(10552.503, 9300.469),(10537.485, 9326.479),(10537.485, 9673.518),(10552.503, 9699.528),(10537.485, 9725.539)), -- tube 344
   345 => ((10585.000, 9274.457),(10600.018, 9300.469),(10585.000, 9326.479),(10585.000, 9673.518),(10600.018, 9699.528),(10585.000, 9725.539)), -- tube 345
   346 => ((10615.035, 9274.457),(10630.053, 9300.469),(10615.035, 9326.479),(10615.035, 9673.518),(10630.053, 9699.528),(10615.035, 9725.539)), -- tube 346
   347 => ((10645.070, 9274.457),(10660.088, 9300.469),(10645.070, 9326.479),(10645.070, 9673.518),(10660.088, 9699.528),(10645.070, 9725.539)), -- tube 347
   348 => ((10675.105, 9274.457),(10690.122, 9300.469),(10675.105, 9326.479),(10675.105, 9673.518),(10690.122, 9699.528),(10675.105, 9725.539)), -- tube 348
   349 => ((10705.140, 9274.457),(10720.157, 9300.469),(10705.140, 9326.479),(10705.140, 9673.518),(10720.157, 9699.528),(10705.140, 9725.539)), -- tube 349
   350 => ((10735.175, 9274.457),(10750.192, 9300.469),(10735.175, 9326.479),(10735.175, 9673.518),(10750.192, 9699.528),(10735.175, 9725.539)), -- tube 350
   351 => ((10765.210, 9274.457),(10780.228, 9300.469),(10765.210, 9326.479),(10765.210, 9673.518),(10780.228, 9699.528),(10765.210, 9725.539)), -- tube 351
   352 => ((10795.245, 9274.457),(10810.263, 9300.469),(10795.245, 9326.479),(10795.245, 9673.518),(10810.263, 9699.528),(10795.245, 9725.539)), -- tube 352
   353 => ((10825.280, 9274.457),(10840.298, 9300.469),(10825.280, 9326.479),(10825.280, 9673.518),(10840.298, 9699.528),(10825.280, 9725.539)), -- tube 353
   354 => ((10855.315, 9274.457),(10870.332, 9300.469),(10855.315, 9326.479),(10855.315, 9673.518),(10870.332, 9699.528),(10855.315, 9725.539)), -- tube 354
   355 => ((10885.350, 9274.457),(10900.367, 9300.469),(10885.350, 9326.479),(10885.350, 9673.518),(10900.367, 9699.528),(10885.350, 9725.539)), -- tube 355
   356 => ((10915.385, 9274.457),(10930.402, 9300.469),(10915.385, 9326.479),(10915.385, 9673.518),(10930.402, 9699.528),(10915.385, 9725.539)), -- tube 356
   357 => ((10945.420, 9274.457),(10960.438, 9300.469),(10945.420, 9326.479),(10945.420, 9673.518),(10960.438, 9699.528),(10945.420, 9725.539)), -- tube 357
   358 => ((10975.455, 9274.457),(10990.473, 9300.469),(10975.455, 9326.479),(10975.455, 9673.518),(10990.473, 9699.528),(10975.455, 9725.539)), -- tube 358
   359 => ((11005.490, 9274.457),(11020.508, 9300.469),(11005.490, 9326.479),(11005.490, 9673.518),(11020.508, 9699.528),(11005.490, 9725.539)), -- tube 359
   360 => ((11035.525, 9274.457),(11050.543, 9300.469),(11035.525, 9326.479),(11035.525, 9673.518),(11050.543, 9699.528),(11035.525, 9725.539)), -- tube 360
   361 => ((11065.560, 9274.457),(11080.577, 9300.469),(11065.560, 9326.479),(11065.560, 9673.518),(11080.577, 9699.528),(11065.560, 9725.539)), -- tube 361
   362 => ((11095.595, 9274.457),(11110.612, 9300.469),(11095.595, 9326.479),(11095.595, 9673.518),(11110.612, 9699.528),(11095.595, 9725.539)), -- tube 362
   363 => ((11125.630, 9274.457),(11140.647, 9300.469),(11125.630, 9326.479),(11125.630, 9673.518),(11140.647, 9699.528),(11125.630, 9725.539)), -- tube 363
   364 => ((11155.665, 9274.457),(11170.683, 9300.469),(11155.665, 9326.479),(11155.665, 9673.518),(11170.683, 9699.528),(11155.665, 9725.539)), -- tube 364
   365 => ((11185.700, 9274.457),(11200.718, 9300.469),(11185.700, 9326.479),(11185.700, 9673.518),(11200.718, 9699.528),(11185.700, 9725.539)), -- tube 365
   366 => ((11215.735, 9274.457),(11230.753, 9300.469),(11215.735, 9326.479),(11215.735, 9673.518),(11230.753, 9699.528),(11215.735, 9725.539)), -- tube 366
   367 => ((11245.770, 9274.457),(11260.787, 9300.469),(11245.770, 9326.479),(11245.770, 9673.518),(11260.787, 9699.528),(11245.770, 9725.539)), -- tube 367
   368 => ((11275.805, 9274.457),(11290.822, 9300.469),(11275.805, 9326.479),(11275.805, 9673.518),(11290.822, 9699.528),(11275.805, 9725.539)), -- tube 368
   369 => ((11305.840, 9274.457),(11320.857, 9300.469),(11305.840, 9326.479),(11305.840, 9673.518),(11320.857, 9699.528),(11305.840, 9725.539)), -- tube 369
   370 => ((11335.875, 9274.457),(11350.893, 9300.469),(11335.875, 9326.479),(11335.875, 9673.518),(11350.893, 9699.528),(11335.875, 9725.539)), -- tube 370
   371 => ((11365.910, 9274.457),(11380.928, 9300.469),(11365.910, 9326.479),(11365.910, 9673.518),(11380.928, 9699.528),(11365.910, 9725.539)), -- tube 371
   372 => ((11395.945, 9274.457),(11410.963, 9300.469),(11395.945, 9326.479),(11395.945, 9673.518),(11410.963, 9699.528),(11395.945, 9725.539)), -- tube 372
   373 => ((11425.980, 9274.457),(11440.997, 9300.469),(11425.980, 9326.479),(11425.980, 9673.518),(11440.997, 9699.528),(11425.980, 9725.539)), -- tube 373
   374 => ((11456.015, 9274.457),(11471.032, 9300.469),(11456.015, 9326.479),(11456.015, 9673.518),(11471.032, 9699.528),(11456.015, 9725.539)), -- tube 374
   375 => ((11486.050, 9274.457),(11501.067, 9300.469),(11486.050, 9326.479),(11486.050, 9673.518),(11501.067, 9699.528),(11486.050, 9725.539)), -- tube 375
   376 => ((11516.085, 9274.457),(11531.103, 9300.469),(11516.085, 9326.479),(11516.085, 9673.518),(11531.103, 9699.528),(11516.085, 9725.539)), -- tube 376
   377 => ((11546.120, 9274.457),(11561.138, 9300.469),(11546.120, 9326.479),(11546.120, 9673.518),(11561.138, 9699.528),(11546.120, 9725.539)), -- tube 377
   378 => ((11576.155, 9274.457),(11591.173, 9300.469),(11576.155, 9326.479),(11576.155, 9673.518),(11591.173, 9699.528),(11576.155, 9725.539)), -- tube 378
   379 => ((11606.190, 9274.457),(11621.207, 9300.469),(11606.190, 9326.479),(11606.190, 9673.518),(11621.207, 9699.528),(11606.190, 9725.539)), -- tube 379
   380 => ((11636.225, 9274.457),(11651.242, 9300.469),(11636.225, 9326.479),(11636.225, 9673.518),(11651.242, 9699.528),(11636.225, 9725.539)), -- tube 380
   381 => ((11666.260, 9274.457),(11681.277, 9300.469),(11666.260, 9326.479),(11666.260, 9673.518),(11681.277, 9699.528),(11666.260, 9725.539)), -- tube 381
   382 => ((11696.295, 9274.457),(11711.312, 9300.469),(11696.295, 9326.479),(11696.295, 9673.518),(11711.312, 9699.528),(11696.295, 9725.539)), -- tube 382
   383 => ((11726.330, 9274.457),(11741.348, 9300.469),(11726.330, 9326.479),(11726.330, 9673.518),(11741.348, 9699.528),(11726.330, 9725.539)), -- tube 383
   384 => ((11756.365, 9274.457),(11771.383, 9300.469),(11756.365, 9326.479),(11756.365, 9673.518),(11771.383, 9699.528),(11756.365, 9725.539)), -- tube 384
   385 => ((11786.400, 9274.457),(11801.418, 9300.469),(11786.400, 9326.479),(11786.400, 9673.518),(11801.418, 9699.528),(11786.400, 9725.539)), -- tube 385
   386 => ((11816.435, 9274.457),(11831.452, 9300.469),(11816.435, 9326.479),(11816.435, 9673.518),(11831.452, 9699.528),(11816.435, 9725.539)), -- tube 386
   387 => ((11846.470, 9274.457),(11861.487, 9300.469),(11846.470, 9326.479),(11846.470, 9673.518),(11861.487, 9699.528),(11846.470, 9725.539)), -- tube 387
   388 => ((11876.505, 9274.457),(11891.522, 9300.469),(11876.505, 9326.479),(11876.505, 9673.518),(11891.522, 9699.528),(11876.505, 9725.539)), -- tube 388
   389 => ((11906.540, 9274.457),(11921.558, 9300.469),(11906.540, 9326.479),(11906.540, 9673.518),(11921.558, 9699.528),(11906.540, 9725.539)), -- tube 389
   390 => ((11936.575, 9274.457),(11951.593, 9300.469),(11936.575, 9326.479),(11936.575, 9673.518),(11951.593, 9699.528),(11936.575, 9725.539)), -- tube 390
   391 => ((11966.610, 9274.457),(11981.628, 9300.469),(11966.610, 9326.479),(11966.610, 9673.518),(11981.628, 9699.528),(11966.610, 9725.539)), -- tube 391
   392 => ((11996.645, 9274.457),(12011.662, 9300.469),(11996.645, 9326.479),(11996.645, 9673.518),(12011.662, 9699.528),(11996.645, 9725.539)), -- tube 392
   393 => ((12026.680, 9274.457),(12041.697, 9300.469),(12026.680, 9326.479),(12026.680, 9673.518),(12041.697, 9699.528),(12026.680, 9725.539)), -- tube 393
   394 => ((12056.715, 9274.457),(12071.732, 9300.469),(12056.715, 9326.479),(12056.715, 9673.518),(12071.732, 9699.528),(12056.715, 9725.539)), -- tube 394
   395 => ((12086.750, 9274.457),(12101.768, 9300.469),(12086.750, 9326.479),(12086.750, 9673.518),(12101.768, 9699.528),(12086.750, 9725.539)), -- tube 395
   396 => ((12116.785, 9274.457),(12131.803, 9300.469),(12116.785, 9326.479),(12116.785, 9673.518),(12131.803, 9699.528),(12116.785, 9725.539)), -- tube 396
   397 => ((12146.820, 9274.457),(12161.838, 9300.469),(12146.820, 9326.479),(12146.820, 9673.518),(12161.838, 9699.528),(12146.820, 9725.539)), -- tube 397
   398 => ((12176.855, 9274.457),(12191.872, 9300.469),(12176.855, 9326.479),(12176.855, 9673.518),(12191.872, 9699.528),(12176.855, 9725.539)), -- tube 398
   399 => ((12206.890, 9274.457),(12221.907, 9300.469),(12206.890, 9326.479),(12206.890, 9673.518),(12221.907, 9699.528),(12206.890, 9725.539))  -- tube 399
  );


 end package TC_B3A_pkg.vhd;
