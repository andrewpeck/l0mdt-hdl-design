module gf_add_3(op1, op2, res);

// -------------------------------------------------------------------------- //
// ------------- Triple Modular Redundancy Generator Directives ------------- //
// -------------------------------------------------------------------------- //
// tmrg do_not_touch
// -------------------------------------------------------------------------- //

	input      [2:0] op1; 
	input      [2:0] op2; 
	output     [2:0] res;

	assign res = op1 ^ op2;

endmodule
