library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.board_pkg_common.all;

package board_pkg is

  constant c_NUM_MGTS                 : integer := 44 + 32;
  constant c_NUM_REFCLKS              : integer := (c_NUM_MGTS/4);

  constant c_MGT_MAP : mgt_inst_array_t (c_NUM_MGTS-1 downto 0) := (

-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    0      => (MGT_LPGBT         , 0      , GTH     , 0 , 0)  ,
    1      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 1)  ,
    2      => (MGT_LPGBT         , 0      , GTH     , 0 , 2)  ,
    3      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 3)  ,
    4      => (MGT_LPGBT         , 1      , GTH     , 0 , 4)  ,
    5      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 5)  ,
    6      => (MGT_LPGBT         , 1      , GTH     , 0 , 6)  ,
    7      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 7)  ,
    8      => (MGT_LPGBT         , 2      , GTH     , 0 , 8)  ,
    9      => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 9)  ,
    10     => (MGT_LPGBT         , 2      , GTH     , 0 , 10) ,
    11     => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 11) ,
    12     => (MGT_LPGBT         , 3      , GTH     , 0 , 12) ,
    13     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 13) ,
    14     => (MGT_LPGBT         , 3      , GTH     , 0 , 14) ,
    15     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 15) ,
    16     => (MGT_LPGBT         , 4      , GTH     , 0 , 16) ,
    17     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 17) ,
    18     => (MGT_LPGBT         , 4      , GTH     , 0 , 18) ,
    19     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 19) ,
    20     => (MGT_LPGBT         , 5      , GTH     , 0 , 20) ,
    21     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 21) ,
    22     => (MGT_LPGBT         , 5      , GTH     , 0 , 22) ,
    23     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 23) ,
    24     => (MGT_LPGBT         , 6      , GTH     , 0 , 24) ,
    25     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 25) ,
    26     => (MGT_LPGBT         , 6      , GTH     , 0 , 26) ,
    27     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 27) ,
    28     => (MGT_LPGBT         , 7      , GTH     , 0 , 28) ,
    29     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 29) ,
    30     => (MGT_LPGBT         , 7      , GTH     , 0 , 30) ,
    31     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 31) ,
    32     => (MGT_SL            , 8      , GTH     , 0 , 32) ,
    33     => (MGT_SL            , 8      , GTH     , 0 , 33) ,
    34     => (MGT_SL            , 8      , GTH     , 0 , 34) ,
    35     => (MGT_SL            , 8      , GTH     , 0 , 35) ,
    36     => (MGT_SL            , 9      , GTH     , 0 , 36) ,
    37     => (MGT_SL            , 9      , GTH     , 0 , 37) ,
    38     => (MGT_SL            , 9      , GTH     , 0 , 38) ,
    39     => (MGT_SL            , 9      , GTH     , 0 , 39) ,
    40     => (MGT_SL            , 10     , GTH     , 0 , 40) ,
    41     => (MGT_SL            , 10     , GTH     , 0 , 41) ,
    42     => (MGT_SL            , 10     , GTH     , 0 , 42) ,
    43     => (MGT_SL            , 10     , GTH     , 0 , 43) ,
-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    44     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 0)  ,
    45     => (MGT_LPGBT         , 11     , GTY     , 0 , 1)  ,
    46     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 2)  ,
    47     => (MGT_LPGBT         , 11     , GTY     , 0 , 3)  ,
    48     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 4)  ,
    49     => (MGT_LPGBT         , 12     , GTY     , 0 , 5)  ,
    50     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 6)  ,
    51     => (MGT_LPGBT         , 12     , GTY     , 0 , 7)  ,
    52     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 8)  ,
    53     => (MGT_LPGBT         , 13     , GTY     , 0 , 9)  ,
    54     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 10) ,
    55     => (MGT_LPGBT         , 13     , GTY     , 0 , 11) ,
    56     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 12) ,
    57     => (MGT_LPGBT         , 14     , GTY     , 0 , 13) ,
    58     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 14) ,
    59     => (MGT_LPGBT         , 14     , GTY     , 0 , 15) ,
    60     => c_mgt_nil ,
    61     => c_mgt_nil ,
    62     => c_mgt_nil ,
    63     => c_mgt_nil ,
    64     => c_mgt_nil ,
    65     => c_mgt_nil ,
    66     => c_mgt_nil ,
    67     => c_mgt_nil ,
    68     => c_mgt_nil ,
    69     => c_mgt_nil ,
    70     => c_mgt_nil ,
    71     => c_mgt_nil ,
    72     => c_mgt_nil ,
    73     => c_mgt_nil ,
    74     => c_mgt_nil ,
    75     => c_mgt_nil ,
    others => c_mgt_nil
    );

  constant c_REFCLK_TYPES : refclk_types_array_t (c_NUM_REFCLKS-1 downto 0) := (
    0      => REFCLK_SYNC320,
    1      => REFCLK_SYNC320,
    2      => REFCLK_SYNC320,
    3      => REFCLK_SYNC320,
    4      => REFCLK_SYNC320,
    others => REFCLK_NIL
    );

  -- FIXME: derive this constant in some sane way
  -- just make it oversized for now and the functions will just ignore the
  -- higher null values... make sure to only specify real things
  constant c_TDC_LINK_MAP : tdc_link_map_array_t (99*14-1 downto 0) := (
    -- TODO: we know that based on the CSM design (once it is final) there are
    -- only certain allowed pairs of even and odd elinks and these can be
    -- derived automatically by just specifying a slot number or something
    --
    -- this is assigned by the global MGT link ID (e.g. 0 to 75 on a ku15p)
    -- mgt link id, even elink #, odd elink #, station
    0      => (link_id => 0, even_elink => 0, odd_elink => 1, station_id => 0),
    1      => (link_id => 0, even_elink => 2, odd_elink => 3, station_id => 0),
    2      => (link_id => 0, even_elink => 4, odd_elink => 5, station_id => 0),
    3      => (link_id => 0, even_elink => 6, odd_elink => 7, station_id => 0),
    4      => (link_id => 0, even_elink => 8, odd_elink => 9, station_id => 0),
    5      => (link_id => 0, even_elink => 10, odd_elink => 11, station_id => 0),
    6      => (link_id => 0, even_elink => 12, odd_elink => 13, station_id => 0),
    7      => (link_id => 0, even_elink => 14, odd_elink => 15, station_id => 0),
    8      => (link_id => 0, even_elink => 16, odd_elink => 17, station_id => 0),
    9      => (link_id => 0, even_elink => 18, odd_elink => 19, station_id => 0),
    10     => (link_id => 0, even_elink => 20, odd_elink => 21, station_id => 0),
    11     => (link_id => 0, even_elink => 22, odd_elink => 23, station_id => 0),
    12     => (link_id => 0, even_elink => 24, odd_elink => 25, station_id => 0),
    13     => (link_id => 0, even_elink => 26, odd_elink => 27, station_id => 0),
    14      => (link_id => 1, even_elink => 0, odd_elink => 1, station_id => 0),
    15      => (link_id => 1, even_elink => 2, odd_elink => 3, station_id => 0),
    16      => (link_id => 1, even_elink => 4, odd_elink => 5, station_id => 0),
    17      => (link_id => 1, even_elink => 6, odd_elink => 7, station_id => 0),
    18      => (link_id => 1, even_elink => 8, odd_elink => 9, station_id => 0),
    19      => (link_id => 1, even_elink => 10, odd_elink => 11, station_id => 0),
    20      => (link_id => 1, even_elink => 12, odd_elink => 13, station_id => 0),
    21      => (link_id => 1, even_elink => 14, odd_elink => 15, station_id => 0),
    22      => (link_id => 1, even_elink => 16, odd_elink => 17, station_id => 0),
    23      => (link_id => 1, even_elink => 18, odd_elink => 19, station_id => 0),
    24     => (link_id => 1, even_elink => 20, odd_elink => 21, station_id => 0),
    25     => (link_id => 1, even_elink => 22, odd_elink => 23, station_id => 0),
    26     => (link_id => 1, even_elink => 24, odd_elink => 25, station_id => 0),
    27     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    28     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    29     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    30     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    31     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    32     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    33     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    34     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    35     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    36     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    37     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    38     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    39     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    40     => (link_id => 2, even_elink => 26, odd_elink => 27, station_id => 0),
    41     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    42     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    43     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    44     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    45     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    46     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    47     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    48     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    49     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    50     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    51     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    52     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    53     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    54     => (link_id => 3, even_elink => 26, odd_elink => 27, station_id => 0),
    55     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    56     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    57     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    58     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    59     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    60     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    61     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    62     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    63     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    64     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    65     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    66     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    67     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    68     => (link_id => 4, even_elink => 26, odd_elink => 27, station_id => 0),
    69     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    70     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    71     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    72     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    73     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    74     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    75     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    76     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    77     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    78     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    79     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    80     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    81     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    82     => (link_id => 5, even_elink => 26, odd_elink => 27, station_id => 0),
    83     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    84     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    85     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    86     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    87     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    88     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    89     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    90     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    91     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    92     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    93     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    94     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    95     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    96     => (link_id => 6, even_elink => 26, odd_elink => 27, station_id => 0),
    97     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    98     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    99     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    100     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    101     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    102     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    103     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    104     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    105     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    106     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    107     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    108     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    109     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    110     => (link_id => 7, even_elink => 26, odd_elink => 27, station_id => 0),
    111     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    112     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    113     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    114     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    115     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    116     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    117     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    118     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    119     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    120     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    121     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    122     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    123     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    124     => (link_id => 8, even_elink => 26, odd_elink => 27, station_id => 0),
    125     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    126     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    127     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    128     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    129     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    130     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    131     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    132     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    133     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    134     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    135     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    136     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    137     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    138     => (link_id => 9, even_elink => 26, odd_elink => 27, station_id => 0),
    139     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    140     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    141     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    142     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    143     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    144     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    145     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    146     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    147     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    148     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    149     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    150     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    151     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    152     => (link_id => 10, even_elink => 26, odd_elink => 27, station_id => 0),
    153     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    154     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    155     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    156     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    157     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    158     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    159     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    160     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    161     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    162     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    163     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    164     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    165     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    166     => (link_id => 11, even_elink => 26, odd_elink => 27, station_id => 0),
    167     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    168     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    169     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    170     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    171     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    172     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    173     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    174     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    175     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    176     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    177     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    178     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    179     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    180     => (link_id => 12, even_elink => 26, odd_elink => 27, station_id => 0),
    181     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    182     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    183     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    184     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    185     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    186     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    187     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    188     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    189     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    190     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    191     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    192     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    193     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    194     => (link_id => 13, even_elink => 26, odd_elink => 27, station_id => 0),
    195     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    196     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    197     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    198     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    199     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    200     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    201     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    202     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    203     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    204     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    205     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    206     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    207     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    208     => (link_id => 14, even_elink => 26, odd_elink => 27, station_id => 0),
    209     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    210     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    211     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    212     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    213     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    214     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    215     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    216     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    217     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    218     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    219     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    220     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    221     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    222     => (link_id => 15, even_elink => 26, odd_elink => 27, station_id => 0),
    223     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    224     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    225     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    226     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    227     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    228     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    229     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    230     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    231     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    232     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    233     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    234     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    235     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    236     => (link_id => 16, even_elink => 26, odd_elink => 27, station_id => 0),
    237     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    238     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    239     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    240     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    241     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    242     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    243     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    244     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    245     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    246     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    247     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    248     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    249     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    250     => (link_id => 17, even_elink => 26, odd_elink => 27, station_id => 0),
    251     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    252     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    253     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    254     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    255     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    256     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    257     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    258     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    259     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    260     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    261     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    262     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    263     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    264     => (link_id => 18, even_elink => 26, odd_elink => 27, station_id => 0),
    265     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    266     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    267     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    268     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    269     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    270     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    271     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    272     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    273     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    274     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    275     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    276     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    277     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    278     => (link_id => 19, even_elink => 26, odd_elink => 27, station_id => 0),
    279     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    280     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    281     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    282     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    283     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    284     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    285     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    286     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    287     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    288     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    289     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    290     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    291     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    292     => (link_id => 20, even_elink => 26, odd_elink => 27, station_id => 0),
    293     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    294     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    295     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    296     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    297     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    298     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    299     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    300     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    301     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    302     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    303     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    304     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    305     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    306     => (link_id => 21, even_elink => 26, odd_elink => 27, station_id => 0),
    307     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    308     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    309     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    310     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    311     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    312     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    313     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    314     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    315     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    316     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    317     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    318     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    319     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    320     => (link_id => 22, even_elink => 26, odd_elink => 27, station_id => 0),
    321     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    322     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    323     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    324     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    325     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    326     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    327     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    328     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    329     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    330     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    331     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    332     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    333     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    334     => (link_id => 23, even_elink => 26, odd_elink => 27, station_id => 0),
    335     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    336     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    337     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    338     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    339     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    340     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    341     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    342     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    343     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    344     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    345     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    346     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    347     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    348     => (link_id => 24, even_elink => 26, odd_elink => 27, station_id => 0),
    349     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    350     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    351     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    352     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    353     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    354     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    355     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    356     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    357     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    358     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    359     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    360     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    361     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    362     => (link_id => 25, even_elink => 26, odd_elink => 27, station_id => 0),
    363     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    364     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    365     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    366     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    367     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    368     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    369     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    370     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    371     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    372     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    373     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    374     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    375     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    376     => (link_id => 26, even_elink => 26, odd_elink => 27, station_id => 0),
    377     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    378     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    379     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    380     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    381     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    382     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    383     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    384     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    385     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    386     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    387     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    388     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    389     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    390     => (link_id => 27, even_elink => 26, odd_elink => 27, station_id => 0),
    391     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    392     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    393     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    394     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    395     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    396     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    397     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    398     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    399     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    400     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    401     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    402     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    403     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    404     => (link_id => 28, even_elink => 26, odd_elink => 27, station_id => 0),
    405     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    406     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    407     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    408     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    409     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    410     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    411     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    412     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    413     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    414     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    415     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    416     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    417     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    418     => (link_id => 29, even_elink => 26, odd_elink => 27, station_id => 0),
    419     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    420     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    421     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    422     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    423     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    424     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    425     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    426     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    427     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    428     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    429     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    430     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    431     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    432     => (link_id => 30, even_elink => 26, odd_elink => 27, station_id => 0),
    433     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    434     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    435     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    436     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    437     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    438     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    439     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    440     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    441     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    442     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    443     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    444     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    445     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),
    446     => (link_id => 31, even_elink => 26, odd_elink => 27, station_id => 0),

    447     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    448     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    449     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    450     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    451     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    452     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    453     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    454     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    455     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    456     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    457     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    458     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    459     => (link_id => 44, even_elink => 26, odd_elink => 27, station_id => 0),
    460     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    461     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    462     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    463     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    464     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    465     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    466     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    467     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    468     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    469     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    470     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    471     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    472     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    473     => (link_id => 45, even_elink => 26, odd_elink => 27, station_id => 0),
    474     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    475     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    476     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    477     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    478     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    479     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    480     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    481     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    482     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    483     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    484     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    485     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    486     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    487     => (link_id => 46, even_elink => 26, odd_elink => 27, station_id => 0),
    488     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    489     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    490     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    491     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    492     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    493     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    494     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    495     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    496     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    497     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    498     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    499     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    500     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    501     => (link_id => 47, even_elink => 26, odd_elink => 27, station_id => 0),
    502     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    503     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    504     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    505     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    506     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    507     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    508     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    509     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    510     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    511     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    512     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    513     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    514     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    515     => (link_id => 48, even_elink => 26, odd_elink => 27, station_id => 0),
    516     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    517     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    518     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    519     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    520     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    521     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    522     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    523     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    524     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    525     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    526     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    527     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    528     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    529     => (link_id => 49, even_elink => 26, odd_elink => 27, station_id => 0),
    530     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    531     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    532     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    533     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    534     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    535     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    536     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    537     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    538     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    539     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    540     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    541     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    542     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    543     => (link_id => 50, even_elink => 26, odd_elink => 27, station_id => 0),
    544     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    545     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    546     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    547     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    548     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    549     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    550     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    551     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    552     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    553     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    554     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    555     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    556     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    557     => (link_id => 51, even_elink => 26, odd_elink => 27, station_id => 0),
    558     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    559     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    560     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    561     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    562     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    563     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    564     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    565     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    566     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    567     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    568     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    569     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    570     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    571     => (link_id => 52, even_elink => 26, odd_elink => 27, station_id => 0),
    572     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    573     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    574     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    575     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    576     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    577     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    578     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    579     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    580     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    581     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    582     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    583     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    584     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    585     => (link_id => 53, even_elink => 26, odd_elink => 27, station_id => 0),
    586     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    587     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    588     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    589     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    590     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    591     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    592     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    593     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    594     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    595     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    596     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    597     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    598     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    599     => (link_id => 54, even_elink => 26, odd_elink => 27, station_id => 0),
    600     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    601     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    602     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    603     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    604     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    605     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    606     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    607     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    608     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    609     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    610     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    611     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    612     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    613     => (link_id => 55, even_elink => 26, odd_elink => 27, station_id => 0),
    614     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    615     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    616     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    617     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    618     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    619     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    620     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    621     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    622     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    623     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    624     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    625     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    626     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    627     => (link_id => 56, even_elink => 26, odd_elink => 27, station_id => 0),
    628     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    629     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    630     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    631     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    632     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    633     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    634     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    635     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    636     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    637     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    638     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    639     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    640     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    641     => (link_id => 57, even_elink => 26, odd_elink => 27, station_id => 0),
    642     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    643     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    644     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    645     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    646     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    647     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    648     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    649     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    650     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    651     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    652     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    653     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    654     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    655     => (link_id => 58, even_elink => 26, odd_elink => 27, station_id => 0),
    656     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    657     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    658     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    659     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    660     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    661     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    662     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    663     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    664     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    665     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    666     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    667     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    668     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    669     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    670     => (link_id => 59, even_elink => 26, odd_elink => 27, station_id => 0),
    others => (-1, -1, -1, -1)
    );

end package board_pkg;
