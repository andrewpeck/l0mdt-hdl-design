../../hal/src/boards/board_pkg_mpi_ku15p.vhd