--------------------------------------------------------------------------------
-- Prototype of functions to convert values to/from text for testbenches
--------------------------------------------------------------------------------
-- original   : Eric Hazen
--      v0.1  : Guillermo   :   added support for TAR
--      v0.2  : Davide      :   CSF version

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;

library shared_lib;
use shared_lib.common_ieee_pkg.all;
use shared_lib.l0mdt_constants_pkg.all;
use shared_lib.l0mdt_dataformats_pkg.all;
use shared_lib.common_constants_pkg.all;
use shared_lib.common_types_pkg.all;
use shared_lib.config_pkg.all;
-- use shared_lib.vhdl2008_functions_pkg.all;
use shared_lib.detector_param_pkg.all;

library project_lib;
use project_lib.gldl_ult_tp_sim_pkg.all;

package csf_textio_pkg is

  procedure READ(L:inout LINE; HIT : out heg2sfhit_rt, SEED : out heg2sfslc_rt, EOF : out std_logic);

  procedure READ(L:inout LINE; VALUE : out input_slc_b_rt);

  -- HEG 2 SF
  procedure WRITEHEADER(L:inout LINE; VALUE : in out_heg_bm_hit_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_hit_sim_rt);

  procedure WRITEHEADER(L:inout LINE; VALUE : in out_heg_bm_slc_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_slc_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_ctrl_sim_rt);
  
  -- PT IN
  procedure WRITEHEADER(L:inout LINE; VALUE : in in_pt_pt2sf_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in in_pt_pt2sf_sim_rt);

  procedure WRITEHEADER(L:inout LINE; VALUE : in in_pt_mpl_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in in_pt_mpl_sim_rt);

  -- MTC IN
  procedure WRITEHEADER(L:inout LINE; VALUE : in in_mtc_pt_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in in_mtc_pt_sim_rt);

  procedure WRITEHEADER(L:inout LINE; VALUE : in in_mtc_mpl_sim_rt);
  procedure WRITE(L:inout LINE; VALUE : in in_mtc_mpl_sim_rt);



end csf_textio_pkg;


package body csf_textio_pkg is

  -----------------------------------------------
  -- read CSF 
  -----------------------------------------------  
  procedure READ(L:inout LINE; HIT : out heg2sfhit_rt, SEED : out heg2sfslc_rt, EOF : out std_logic) is

    variable hit_dv : integer;
    variable hit_ml : integer;
    variable hit_x  : integer;
    variable hit_y  : integer;
    variable hit_r  : integer;
    variable slc_dv : integer;
    variable slc_chamber_id : integer;
    variable slc_chamber_ieta : integer;
    variable slc_vec_pos : integer;
    variable slc_vec_ang : integer;
    variable slc_hewindow_pos : integer;
    variable eof : integer;

    variable mdt_ToA  : integer;
    -- variable tdc_time     : integer;
    -- variable space        : string(8 downto 1);
    -- variable c_Station    : string(1 downto 1);
    variable i_station        : integer;
    variable Chamber_id       : integer;
    variable Chamber_ieta     : integer;
    variable mdt_time_coarse  : integer;
    variable mdt_time_fine    : integer;
    variable tube_global      : integer;
    variable tube_local       : integer;
    variable tube_layer       : integer;
    variable tube_z           : integer;
    variable tube_rho         : integer;
    variable drift_time       : real;
    variable event            : integer;
    variable muonFixedId      : integer;
    variable csm              : integer;
    variable mezz             : integer;
    variable channel          : integer;
    variable t0               : real;
    variable TOF              : real;

    variable dummy_text  : string(1 to 100);
    variable ok : boolean;

    -- variable
  begin
    -- Event
    -- READ(L, event);
    -- Hit Data Valid
    READ(L, hit_dv);
    -- Hit Multilayer
    READ(L, hit_ml);
    -- Hit Local X
    READ(L, hit_x);
    -- Hit Local Y
    READ(L, hit_y);
    -- Hit Radius
    READ(L, hit_r);
    -- SLC dv
    READ(L, slc_dv);
    -- ChamberId < Chamber ID using L0MDT numbering scheme
    READ(L, slc_chamber_id);
    -- Chamber_iEta < iEta index of the chamber [0,7]. Based on 1st layer of tube.
    READ(L, slc_chamber_ieta);
    -- SLC vec_pos
    READ(L, slc_vec_pos);
    -- SLC vec_ang (mbar for csf)
    READ(L, slc_vec_ang);
    -- SLC HE window pos
    READ(L, slc_hewindow_pos);
    -- EOF
    READ(L, file_eof);
    
    HIT := (
      data_valid => std_logic(to_unsigned(hit_dv,1)),
      mlayer => std_logic(to_unsigned(hit_ml,1)),
      localx => to_unsigned(hit_x, HEG2SFHIT_LOCALX_LEN),
      localy => to_unsigned(hit_y, HEG2SFHIT_LOCALY_LEN),
      radius => to_unsigned(hit_r, HEG2SFHIT_RADIUS_LEN)
    )

    SEED := (
      data_valid => std_logic(to_unsigned(slc_dv,1)),
      mdtid => (
        chamber_id => to_unsigned(slc_chamber_id, VEC_MDTID_CHAMBER_ID_LEN),
        chamber_ieta => to_unsigned(slc_chamber_ieta, VEC_MDTID_CHAMBER_IETA_LEN)
        ),
      vec_pos => to_unsigned(slc_vec_pos, UCM2HPS_VEC_POS_LEN),
      vec_ang => to_unsigned(slc_vec_ang, UCM2HPS_VEC_ANG_LEN),
      hewindow_pos => to_unsigned(slc_hewindow_pos, HEG2SFSLC_HEWINDOW_POS_LEN)
    )

    EOF := std_logic(to_unsigned(file_eof, 1));

  end procedure;

  -----------------------------------------------
  -- read SLC 
  -----------------------------------------------  
  procedure READ(L:inout LINE; VALUE : out input_slc_b_rt) is
    variable BCID         : integer; 
    variable ToA          : integer; 
    variable nTC          : integer; 
    variable TC_sent      : integer; 
    variable TC_id        : integer; 
    variable Eta          : real; 
    variable Phi          : real; 
    variable pT_thr       : integer; 
    variable Charge       : integer; 
    variable Coincidence  : integer; 
    variable z_RPC0       : integer; 
    variable z_RPC1       : integer; 
    variable z_RPC2       : integer; 
    variable z_RPC3       : integer; 

    variable header       : sl_header_rt;
    variable trailer      : sl_trailer_rt;
    variable common       : slc_common_rt;
    variable specific     : slc_barrel_rt;
    
    variable tcoverflow : std_logic;


  begin
    READ( L , BCID );
    READ( L , ToA );
    READ( L , nTC );
    READ( L , TC_sent );
    READ( L , TC_id );
    READ( L , Eta );
    READ( L , Phi );
    READ( L , pT_thr );
    READ( L , Charge );
    READ( L , Coincidence );
    READ( L , z_RPC0 );
    READ( L , z_RPC1 );
    READ( L , z_RPC2 );
    READ( L , z_RPC3 );

    if nTC > 3 then 
      tcoverflow := '1';
    else
      tcoverflow := '0';
    end if;

    header := (
      h_reserved => (others => '1'),
      tcoverflow => tcoverflow,
      nmtc_sl    => to_unsigned(nTC, SL_HEADER_NSLC_LEN),
      nmtc_mdt   => (others => '1'),
      nslc       => (others => '1'),
      bcid       => to_unsigned(BCID, SL_HEADER_BCID_LEN)
    );

    trailer :=(
      t_reserved => (others => '1'),
      crc        => (others => '1'),
      fiberid    => (others => '1'),
      slid       => (others => '1'),
      comma      => (others => '1')
    );

    common := (
      header      => header,
      slcid       => to_unsigned(TC_id, SL_HEADER_NSLC_LEN),
      tcsent      => std_logic(to_unsigned(TC_sent,1)(0)),
      poseta      => to_signed(integer(Eta * SLC_COMMON_POSETA_MULT), SLC_COMMON_POSETA_LEN) ,
      posphi      => to_unsigned(integer((Phi * SLC_COMMON_POSPHI_MULT/1000.0)), SLC_COMMON_POSPHI_LEN) , 
      sl_pt       => ( others => '0'),
      sl_ptthresh => to_unsigned(pT_thr, SLC_COMMON_SL_PTTHRESH_LEN) , 
      sl_charge   => std_logic(to_unsigned(Charge,1)(0)), 
      cointype    => std_logic_vector(to_unsigned(Coincidence,SLC_COMMON_COINTYPE_LEN)), 
      trailer     => trailer
    );

    specific :=(
      -- b_reserved  => (others => '0'),
      rpc0_posz   => to_signed(integer(real(z_RPC0) * SLC_Z_RPC_MULT) ,SLC_BARREL_RPC0_POSZ_LEN) ,
      rpc1_posz   => to_signed(integer(real(z_RPC1) * SLC_Z_RPC_MULT) ,SLC_BARREL_RPC1_POSZ_LEN) ,
      rpc2_posz   => to_signed(integer(real(z_RPC2) * SLC_Z_RPC_MULT) ,SLC_BARREL_RPC2_POSZ_LEN) ,
      rpc3_posz   => to_signed(integer(real(z_RPC3) * SLC_Z_RPC_MULT) ,SLC_BARREL_RPC3_POSZ_LEN)
    );

    VALUE := (
      ToA => to_unsigned(ToA , 64) , 
      slc => (
        data_Valid  => '1',
        common      => common,
        specific    => std_logic_vector(vectorify(specific))
      )
    );

    report "##### SLC : " & integer'image(BCID) &
    " - " & integer'image(ToA) &
    " - " & integer'image(nTC) &
    " - " & integer'image(TC_sent) &
    " - " & integer'image(TC_id) &
    " - " & real'image(Eta) &
    " - " & real'image(Phi) &
    " - " & integer'image(pT_thr) &
    " - " & integer'image(Charge) &
    " - " & integer'image(Coincidence) &
    " - " & integer'image(z_RPC0) &
    " - " & integer'image(z_RPC1) &
    " - " & integer'image(z_RPC2) &
    " - " & integer'image(z_RPC3);
  end procedure;
  -----------------------------------------------
  -- HEG(HIT) 2 SF
  -----------------------------------------------  
  procedure WRITEHEADER(L:inout LINE; VALUE : in out_heg_bm_hit_sim_rt) is
  begin
    -- SWRITE(L, "#");
    -- SWRITE(L, "FLAG");
    SWRITE(L, "ToA");
    WRITE(L, ',');
    SWRITE(L, "station");
    WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "data_valid");
    WRITE(L, ',');
    SWRITE(L, "mlayer");
    WRITE(L, ',');
    SWRITE(L, "localx");
    WRITE(L, ',');
    SWRITE(L, "localy");
    WRITE(L, ',');
    SWRITE(L, "radius");
  end procedure;
  
  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_hit_sim_rt) is

    variable ToA      : unsigned(64-1 downto 0);
    variable station  : unsigned(4-1 downto 0);
    variable thread   : unsigned(4-1 downto 0);
    variable mlayer   : std_logic;
    variable localx   : unsigned(HEG2SFHIT_LOCALX_LEN-1 downto 0);
    variable localy   : unsigned(HEG2SFHIT_LOCALY_LEN-1 downto 0);
    variable radius   : unsigned(HEG2SFHIT_RADIUS_LEN-1 downto 0);
    variable data_valid : std_logic;

  begin

    ToA     := VALUE.ToA;
    station := VALUE.station;
    thread  := VALUE.thread;
    data_valid  := VALUE.data.data_valid;
    mlayer  := VALUE.data.mlayer;
    localx  := VALUE.data.localx;
    localy  := VALUE.data.localy;
    radius  := VALUE.data.radius;

    -- SWRITE(L, " HIT: ");
    -- SWRITE(L, "NONE");
    WRITE(L, to_integer( ToA));
    WRITE(L, ',');
    WRITE(L, to_integer( station));
    WRITE(L, ',');
    WRITE(L, to_integer( thread));
    WRITE(L, ',');
    WRITE(L, data_valid);
    WRITE(L, ',');
    WRITE(L, mlayer);
    WRITE(L, ',');
    WRITE(L, to_integer( localx));
    WRITE(L, ',');
    WRITE(L, to_integer( localy));
    WRITE(L, ',');
    WRITE(L, to_integer( radius));

  end procedure;
  -----------------------------------------------
  -- HEG(SLC) 2 SF 
  -----------------------------------------------  
  procedure WRITEHEADER(L:inout LINE; VALUE : in out_heg_bm_slc_sim_rt) is
  begin

    SWRITE(L, "ToA");
    WRITE(L, ',');
    SWRITE(L, "FLAG");
    WRITE(L, ',');

    SWRITE(L, "station");
    WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "slcid");
    WRITE(L, ',');
    SWRITE(L, "slid");
    WRITE(L, ',');
    SWRITE(L, "bcid");
    WRITE(L, ',');
    SWRITE(L, "mdtseg_dest");
    WRITE(L, ',');
    SWRITE(L, "chamber_id");
    WRITE(L, ',');
    SWRITE(L, "chamber_ieta");
    WRITE(L, ',');
    SWRITE(L, "vec_pos");
    WRITE(L, ',');
    SWRITE(L, "vec_ang");
    WRITE(L, ',');
    SWRITE(L, "hewindow_pos");
  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_slc_sim_rt) is

    variable ToA          : unsigned(64-1 downto 0);
    variable station      : unsigned(4-1 downto 0);
    variable thread       : unsigned(4-1 downto 0);
    variable slcid        : unsigned(SLC_COMMON_SLCID_LEN-1 downto 0);
    variable slid         : unsigned(SL_TRAILER_SLID_LEN-1 downto 0);
    variable bcid         : unsigned(SL_HEADER_BCID_LEN-1 downto 0);
    variable mdtseg_dest  : std_logic_vector(HEG2SFSLC_MDTSEG_DEST_LEN-1 downto 0);
    variable chamber_id   : unsigned(VEC_MDTID_CHAMBER_ID_LEN-1 downto 0);
    variable chamber_ieta : unsigned(VEC_MDTID_CHAMBER_IETA_LEN-1 downto 0);
    variable vec_pos      : unsigned(UCM2HPS_VEC_POS_LEN-1 downto 0);
    variable vec_ang      : unsigned(UCM2HPS_VEC_ANG_LEN-1 downto 0);
    variable hewindow_pos : unsigned(HEG2SFSLC_HEWINDOW_POS_LEN-1 downto 0);

  begin

    ToA           := VALUE.ToA;
    station       := VALUE.station;
    thread        := VALUE.thread;
    slcid         := VALUE.data.muid.slcid;
    slid          := VALUE.data.muid.slid;
    bcid          := VALUE.data.muid.bcid;
    mdtseg_dest   := VALUE.data.mdtseg_dest; 
    chamber_id    := VALUE.data.mdtid.chamber_id;
    chamber_ieta  := VALUE.data.mdtid.chamber_ieta;
    vec_pos       := VALUE.data.vec_pos;
    vec_ang       := VALUE.data.vec_ang;
    hewindow_pos  := VALUE.data.hewindow_pos;

    WRITE(L, to_integer( ToA));
    WRITE(L, ',');
    SWRITE(L, "SOF");
    WRITE(L, ',');
    WRITE(L, to_integer( station));
    WRITE(L, ',');
    WRITE(L, to_integer( thread));
    WRITE(L, ',');
    WRITE(L, to_integer( slcid));
    WRITE(L, ',');
    WRITE(L, to_integer( slid));
    WRITE(L, ',');
    WRITE(L, to_integer( bcid));
    WRITE(L, ',');
    WRITE(L, to_integer(unsigned(mdtseg_dest)));
    WRITE(L, ',');
    WRITE(L, to_integer( chamber_id));
    WRITE(L, ',');
    WRITE(L, to_integer( chamber_ieta));
    WRITE(L, ',');
    WRITE(L, to_integer( vec_pos));
    WRITE(L, ',');
    WRITE(L, to_integer( vec_ang));
    WRITE(L, ',');
    WRITE(L, to_integer( hewindow_pos));

  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in out_heg_bm_ctrl_sim_rt) is

    variable ToA          : unsigned(64-1 downto 0);
    variable station      : unsigned(4-1 downto 0);
    variable thread       : unsigned(4-1 downto 0);
    variable slcid        : unsigned(SLC_COMMON_SLCID_LEN-1 downto 0);
    variable slid         : unsigned(SL_TRAILER_SLID_LEN-1 downto 0);
    variable bcid         : unsigned(SL_HEADER_BCID_LEN-1 downto 0);
    variable mdtseg_dest  : std_logic_vector(HEG2SFSLC_MDTSEG_DEST_LEN-1 downto 0);
    variable chamber_id   : unsigned(VEC_MDTID_CHAMBER_ID_LEN-1 downto 0);
    variable chamber_ieta : unsigned(VEC_MDTID_CHAMBER_IETA_LEN-1 downto 0);
    variable vec_pos      : unsigned(UCM2HPS_VEC_POS_LEN-1 downto 0);
    variable vec_ang      : unsigned(UCM2HPS_VEC_ANG_LEN-1 downto 0);
    variable hewindow_pos : unsigned(HEG2SFSLC_HEWINDOW_POS_LEN-1 downto 0);

  begin

    ToA           := VALUE.ToA;
    station       := VALUE.station;
    thread        := VALUE.thread;
    slcid         := VALUE.data.muid.slcid;
    slid          := VALUE.data.muid.slid;
    bcid          := VALUE.data.muid.bcid;
    mdtseg_dest   := VALUE.data.mdtseg_dest; 
    chamber_id    := VALUE.data.mdtid.chamber_id;
    chamber_ieta  := VALUE.data.mdtid.chamber_ieta;
    vec_pos       := VALUE.data.vec_pos;
    vec_ang       := VALUE.data.vec_ang;
    hewindow_pos  := VALUE.data.hewindow_pos;

    WRITE(L, to_integer( ToA));
    WRITE(L, ',');
    SWRITE(L, "EOF");
    WRITE(L, ',');
    WRITE(L, to_integer( station));
    WRITE(L, ',');
    WRITE(L, to_integer( thread));
    WRITE(L, ',');
    WRITE(L, to_integer( slcid));
    WRITE(L, ',');
    WRITE(L, to_integer( slid));
    WRITE(L, ',');
    WRITE(L, to_integer( bcid));
    WRITE(L, ',');
    WRITE(L, to_integer(unsigned(mdtseg_dest)));
    WRITE(L, ',');
    WRITE(L, to_integer( chamber_id));
    WRITE(L, ',');
    WRITE(L, to_integer( chamber_ieta));
    WRITE(L, ',');
    WRITE(L, to_integer( vec_pos));
    WRITE(L, ',');
    WRITE(L, to_integer( vec_ang));
    WRITE(L, ',');
    WRITE(L, to_integer( hewindow_pos));

  end procedure;

  -----------------------------------------------
  -- SF 2 PT 
  -----------------------------------------------  


  procedure WRITEHEADER(L:inout LINE; VALUE : in in_pt_pt2sf_sim_rt) is
  begin

    -- SWRITE(L, "# ");
    -- SWRITE(L, "FLAG");
    -- WRITE(L, ',');
    SWRITE(L, "ToA");
    WRITE(L, ',');
    SWRITE(L, "station");
    WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "slcid");
    WRITE(L, ',');
    SWRITE(L, "slid");
    WRITE(L, ',');
    SWRITE(L, "bcid");
    -- WRITE(L, ',');
    -- SWRITE(L, "mdtseg_dest");
    WRITE(L, ',');
    SWRITE(L, "chamber_id");
    WRITE(L, ',');
    SWRITE(L, "chamber_ieta");
    WRITE(L, ',');
    SWRITE(L, "segpos");
    WRITE(L, ',');
    SWRITE(L, "segangle");
    WRITE(L, ',');
    SWRITE(L, "segquality");
  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in in_pt_pt2sf_sim_rt) is

    variable ToA          : unsigned(64-1 downto 0);
    variable station      : unsigned(4-1 downto 0);
    variable thread       : unsigned(4-1 downto 0);
    variable slcid        : unsigned(SLC_COMMON_SLCID_LEN-1 downto 0);
    variable slid         : unsigned(SL_TRAILER_SLID_LEN-1 downto 0);
    variable bcid         : unsigned(SL_HEADER_BCID_LEN-1 downto 0);
    -- variable mdtseg_dest  : std_logic_vector(HEG2SFSLC_MDTSEG_DEST_LEN-1 downto 0);
    variable chamber_id   : unsigned(VEC_MDTID_CHAMBER_ID_LEN-1 downto 0);
    variable chamber_ieta : unsigned(VEC_MDTID_CHAMBER_IETA_LEN-1 downto 0);
    -- variable vec_pos      : unsigned(UCM2HPS_VEC_POS_LEN-1 downto 0);
    -- variable vec_ang      : unsigned(UCM2HPS_VEC_ANG_LEN-1 downto 0);
    -- variable hewindow_pos : unsigned(HEG2SFSLC_HEWINDOW_POS_LEN-1 downto 0);
    variable segpos       : unsigned(SF2PTCALC_SEGPOS_LEN-1 downto 0);
    variable segangle     : unsigned(SF2PTCALC_SEGANGLE_LEN-1 downto 0);
    variable segquality   : std_logic;

  begin

    ToA           := VALUE.ToA;
    station       := VALUE.station;
    thread        := VALUE.thread;
    slcid         := VALUE.data.muid.slcid;
    slid          := VALUE.data.muid.slid;
    bcid          := VALUE.data.muid.bcid;
    -- mdtseg_dest   := VALUE.data.mdtseg_dest; 
    chamber_id    := VALUE.data.mdtid.chamber_id;
    chamber_ieta  := VALUE.data.mdtid.chamber_ieta;
    segpos        := VALUE.data.segpos;
    segangle      := VALUE.data.segangle;
    segquality    := VALUE.data.segquality;


    WRITE(L, to_integer( ToA));
    WRITE(L, ',');
    WRITE(L, to_integer( station));
    WRITE(L, ',');
    WRITE(L, to_integer( thread));
    WRITE(L, ',');
    WRITE(L, to_integer( slcid));
    WRITE(L, ',');
    WRITE(L, to_integer( slid));
    WRITE(L, ',');
    WRITE(L, to_integer( bcid));
    WRITE(L, ',');
    -- WRITE(L, to_integer(unsigned(mdtseg_dest)));
    -- WRITE(L, ',');
    WRITE(L, to_integer( chamber_id));
    WRITE(L, ',');
    WRITE(L, to_integer( chamber_ieta));
    WRITE(L, ',');
    WRITE(L, to_integer( segpos));
    WRITE(L, ',');
    WRITE(L, to_integer( segangle));
    WRITE(L, ',');
    WRITE(L, segquality);

  end procedure;

  -----------------------------------------------
  -- MPL 2 PT 
  -----------------------------------------------  

  procedure WRITEHEADER(L:inout LINE; VALUE : in in_pt_mpl_sim_rt) is
  begin

    -- SWRITE(L, "# ");
    -- SWRITE(L, "FLAG");
    -- WRITE(L, ',');
    SWRITE(L, "ToA");
    WRITE(L, ',');
    -- SWRITE(L, "station");
    -- WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "slcid");
    WRITE(L, ',');
    SWRITE(L, "slid");
    WRITE(L, ',');
    SWRITE(L, "bcid");
    WRITE(L, ',');
    -- SWRITE(L, "mdtseg_dest");
    -- WRITE(L, ',');
    SWRITE(L, "phimod");
    WRITE(L, ',');
    SWRITE(L, "sl_charge");
    WRITE(L, ',');
    SWRITE(L, "nswseg_poseta");
    WRITE(L, ',');
    SWRITE(L, "nswseg_posphi");
    WRITE(L, ',');
    SWRITE(L, "nswseg_angdtheta");
  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in in_pt_mpl_sim_rt) is

    variable ToA              : unsigned(64-1 downto 0);
    variable station          : unsigned(4-1 downto 0);
    variable thread           : unsigned(4-1 downto 0);
    -- variable busy             : std_logic;
    -- variable process_ch       : std_logic_vector(UCM2PL_PROCESS_CH_LEN-1 downto 0);
    variable slcid            : unsigned(SLC_COMMON_SLCID_LEN-1 downto 0);
    variable slid             : unsigned(SL_TRAILER_SLID_LEN-1 downto 0);
    variable bcid             : unsigned(SL_HEADER_BCID_LEN-1 downto 0);
    variable phimod           : signed(UCM2PL_PHIMOD_LEN-1 downto 0);
    variable sl_charge        : std_logic;
    variable nswseg_poseta    : unsigned(SLC_ENDCAP_NSWSEG_POSETA_LEN-1 downto 0);
    variable nswseg_posphi    : unsigned(SLC_ENDCAP_NSWSEG_POSPHI_LEN-1 downto 0);
    variable nswseg_angdtheta : signed(SLC_ENDCAP_NSWSEG_ANGDTHETA_LEN-1 downto 0);
  

  begin

    ToA               := VALUE.ToA;
    -- station           := VALUE.station;
    thread            := VALUE.thread;
    -- busy          := VALUE.data.busy;
    -- process_ch    := VALUE.data.process_ch;
    slcid             := VALUE.data.muid.slcid;
    slid              := VALUE.data.muid.slid;
    bcid              := VALUE.data.muid.bcid;
    phimod            := VALUE.data.phimod; 
    sl_charge         := VALUE.data.sl_charge;
    nswseg_poseta     := VALUE.data.nswseg_poseta;
    nswseg_posphi     := VALUE.data.nswseg_posphi;
    nswseg_angdtheta  := VALUE.data.nswseg_angdtheta;

    WRITE(L, to_integer( ToA));
    WRITE(L, ',');
    -- WRITE(L, to_integer( station));
    -- WRITE(L, ',');
    WRITE(L, to_integer( thread));
    WRITE(L, ',');
    -- WRITE(L, to_integer( slcid));
    -- WRITE(L, ',');
    -- WRITE(L, to_integer( slcid));
    -- WRITE(L, ',');
    WRITE(L, to_integer( slcid));
    WRITE(L, ',');
    WRITE(L, to_integer( slid));
    WRITE(L, ',');
    WRITE(L, to_integer( bcid));
    WRITE(L, ',');
    -- WRITE(L, to_integer(unsigned(mdtseg_dest)));
    -- WRITE(L, ',');
    WRITE(L, to_integer( phimod));
    WRITE(L, ',');
    WRITE(L, sl_charge);
    WRITE(L, ',');
    WRITE(L, to_integer( nswseg_poseta));
    WRITE(L, ',');
    WRITE(L, to_integer( nswseg_posphi));
    WRITE(L, ',');
    WRITE(L, to_integer( nswseg_angdtheta));

  end procedure;
  -----------------------------------------------
  -- PT 2 MTCB
  -----------------------------------------------  
  procedure WRITEHEADER(L:inout LINE; VALUE : in in_mtc_pt_sim_rt) is
  begin

    SWRITE(L, "ToA");
    WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "slcid");
    WRITE(L, ',');
    SWRITE(L, "slid");
    WRITE(L, ',');
    SWRITE(L, "bcid");
    WRITE(L, ',');
    SWRITE(L, "mdt_eta");
    WRITE(L, ',');
    SWRITE(L, "mdt_pt");
    WRITE(L, ',');
    SWRITE(L, "mdt_ptthresh");
    WRITE(L, ',');
    SWRITE(L, "mdt_charge");
    WRITE(L, ',');
    SWRITE(L, "mdt_nsegments");
    WRITE(L, ',');
    SWRITE(L, "mdt_quality");

  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in in_mtc_pt_sim_rt) is


  begin

    WRITE(L, to_integer( VALUE.ToA));
    WRITE(L, ',');
    WRITE(L, to_integer( VALUE.thread));
    WRITE(L, ',');
    WRITE(L, VALUE.data.muid.slcid);
    WRITE(L, ',');      
    WRITE(L, VALUE.data.muid.slid);
    WRITE(L, ',');      
    WRITE(L, VALUE.data.muid.bcid);
    WRITE(L, ',');    
    WRITE(L, to_integer( VALUE.data.mdt_eta));
    WRITE(L, ',');
    WRITE(L, to_integer( VALUE.data.mdt_pt));
    WRITE(L, ',');
    WRITE(L, to_integer( VALUE.data.mdt_ptthresh));
    WRITE(L, ',');
    WRITE(L, VALUE.data.mdt_charge);
    WRITE(L, ',');
    WRITE(L, to_integer( VALUE.data.mdt_nsegments));
    WRITE(L, ',');
    WRITE(L, to_integer( unsigned(VALUE.data.mdt_quality)));

  end procedure;
  -----------------------------------------------
  -- MPL 2 MTCB
  -----------------------------------------------  
  procedure WRITEHEADER(L:inout LINE; VALUE : in in_mtc_mpl_sim_rt) is
  begin

    SWRITE(L, "ToA");
    WRITE(L, ',');
    SWRITE(L, "thread");
    WRITE(L, ',');
    SWRITE(L, "processed");
    WRITE(L, ',');
    SWRITE(L, "tcoverflow");
    WRITE(L, ',');
    SWRITE(L, "nmtc_sl");
    WRITE(L, ',');
    SWRITE(L, "nmtc_mdt");
    WRITE(L, ',');
    SWRITE(L, "nslc");
    WRITE(L, ',');
    SWRITE(L, "bcid");
    WRITE(L, ',');
    SWRITE(L, "slcid");
    WRITE(L, ',');
    SWRITE(L, "tcsent");
    WRITE(L, ',');
    SWRITE(L, "poseta");
    WRITE(L, ',');
    SWRITE(L, "posphi");
    WRITE(L, ',');
    SWRITE(L, "sl_pt");
    WRITE(L, ',');
    SWRITE(L, "sl_ptthresh");
    WRITE(L, ',');
    SWRITE(L, "sl_charge");
    WRITE(L, ',');
    SWRITE(L, "cointype");

  end procedure;

  procedure WRITE(L:inout LINE; VALUE : in in_mtc_mpl_sim_rt) is
    -- variable ToA              : unsigned(64-1 downto 0);
    -- variable station          : unsigned(4-1 downto 0);
    -- variable thread           : unsigned(4-1 downto 0);

    variable slc_common_r     : slc_common_rt;
    variable sl_header_r      : sl_header_rt;

  begin

    slc_common_r  := VALUE.data.common;
    sl_header_r   := slc_common_r.header;

    WRITE(L, to_integer( VALUE.ToA));
    WRITE(L, ',');
    WRITE(L, to_integer( VALUE.thread));
    WRITE(L, ',');
    WRITE(L, VALUE.data.busy);
    WRITE(L, ',');    
    WRITE(L, to_integer( unsigned( VALUE.data.process_ch)));
    WRITE(L, ',');

    WRITE(L, sl_header_r.tcoverflow);
    WRITE(L, ',');
    WRITE(L, to_integer( unsigned(sl_header_r.nmtc_sl)));
    WRITE(L, ',');
    WRITE(L, to_integer( unsigned(sl_header_r.nmtc_mdt)));
    WRITE(L, ',');
    WRITE(L, to_integer( unsigned(sl_header_r.nslc)));
    WRITE(L, ',');
    WRITE(L, to_integer( unsigned(sl_header_r.bcid)));
    WRITE(L, ',');

    WRITE(L, to_integer( slc_common_r.slcid));
    WRITE(L, ',');
    WRITE(L, slc_common_r.tcsent);
    WRITE(L, ',');
    WRITE(L, to_integer( slc_common_r.poseta));
    WRITE(L, ',');
    WRITE(L, to_integer( slc_common_r.posphi));
    WRITE(L, ',');
    WRITE(L, to_integer(unsigned(slc_common_r.sl_pt)));
    WRITE(L, ',');    
    WRITE(L, to_integer(unsigned(slc_common_r.sl_ptthresh)));
    WRITE(L, ',');
    WRITE(L, slc_common_r.sl_charge );
    WRITE(L, ',');
    WRITE(L, to_integer(unsigned(slc_common_r.cointype)));

  end procedure;


end gldl_l0mdt_textio_pkg;