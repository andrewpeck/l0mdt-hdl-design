../../hw/tdc/tdc_decoder_wrapper.vhd