library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.board_pkg_common.all;

package board_pkg is

  constant c_NUM_MGTS                 : integer := 44 + 32;
  constant c_NUM_REFCLKS              : integer := (c_NUM_MGTS/4);

  constant c_MGT_MAP : mgt_inst_array_t (c_NUM_MGTS-1 downto 0) := (

-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    0      => (MGT_LPGBT         , 0      , GTH     , 0 , 0)  ,
    1      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 1)  ,
    2      => (MGT_LPGBT         , 0      , GTH     , 0 , 2)  ,
    3      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 3)  ,
    4      => (MGT_LPGBT         , 1      , GTH     , 0 , 4)  ,
    5      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 5)  ,
    6      => (MGT_LPGBT         , 1      , GTH     , 0 , 6)  ,
    7      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 7)  ,
    8      => (MGT_LPGBT         , 2      , GTH     , 0 , 8)  ,
    9      => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 9)  ,
    10     => (MGT_LPGBT         , 2      , GTH     , 0 , 10) ,
    11     => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 11) ,
    12     => (MGT_LPGBT         , 3      , GTH     , 0 , 12) ,
    13     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 13) ,
    14     => (MGT_LPGBT         , 3      , GTH     , 0 , 14) ,
    15     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 15) ,
    16     => (MGT_LPGBT         , 4      , GTH     , 0 , 16) ,
    17     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 17) ,
    18     => (MGT_LPGBT         , 4      , GTH     , 0 , 18) ,
    19     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 19) ,
    20     => (MGT_LPGBT         , 5      , GTH     , 0 , 20) ,
    21     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 21) ,
    22     => (MGT_LPGBT         , 5      , GTH     , 0 , 22) ,
    23     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 23) ,
    24     => (MGT_LPGBT         , 6      , GTH     , 0 , 24) ,
    25     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 25) ,
    26     => (MGT_LPGBT         , 6      , GTH     , 0 , 26) ,
    27     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 27) ,
    28     => (MGT_LPGBT         , 7      , GTH     , 0 , 28) ,
    29     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 29) ,
    30     => (MGT_LPGBT         , 7      , GTH     , 0 , 30) ,
    31     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 31) ,
    32     => (MGT_SL            , 8      , GTH     , 0 , 32) ,
    33     => (MGT_SL            , 8      , GTH     , 0 , 33) ,
    34     => (MGT_SL            , 8      , GTH     , 0 , 34) ,
    35     => (MGT_SL            , 8      , GTH     , 0 , 35) ,
    36     => (MGT_SL            , 9      , GTH     , 0 , 36) ,
    37     => (MGT_SL            , 9      , GTH     , 0 , 37) ,
    38     => (MGT_SL            , 9      , GTH     , 0 , 38) ,
    39     => (MGT_SL            , 9      , GTH     , 0 , 39) ,
    40     => (MGT_SL            , 10     , GTH     , 0 , 40) ,
    41     => (MGT_SL            , 10     , GTH     , 0 , 41) ,
    42     => (MGT_SL            , 10     , GTH     , 0 , 42) ,
    43     => (MGT_SL            , 10     , GTH     , 0 , 43) ,
-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    44     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 0)  ,
    45     => (MGT_LPGBT         , 11     , GTY     , 0 , 1)  ,
    46     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 2)  ,
    47     => (MGT_LPGBT         , 11     , GTY     , 0 , 3)  ,
    48     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 4)  ,
    49     => (MGT_LPGBT         , 12     , GTY     , 0 , 5)  ,
    50     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 6)  ,
    51     => (MGT_LPGBT         , 12     , GTY     , 0 , 7)  ,
    52     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 8)  ,
    53     => (MGT_LPGBT         , 13     , GTY     , 0 , 9)  ,
    54     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 10) ,
    55     => (MGT_LPGBT         , 13     , GTY     , 0 , 11) ,
    56     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 12) ,
    57     => (MGT_LPGBT         , 14     , GTY     , 0 , 13) ,
    58     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 14) ,
    59     => (MGT_LPGBT         , 14     , GTY     , 0 , 15) ,
    60     => c_mgt_nil ,
    61     => c_mgt_nil ,
    62     => c_mgt_nil ,
    63     => c_mgt_nil ,
    64     => c_mgt_nil ,
    65     => c_mgt_nil ,
    66     => c_mgt_nil ,
    67     => c_mgt_nil ,
    68     => c_mgt_nil ,
    69     => c_mgt_nil ,
    70     => c_mgt_nil ,
    71     => c_mgt_nil ,
    72     => c_mgt_nil ,
    73     => c_mgt_nil ,
    74     => c_mgt_nil ,
    75     => c_mgt_nil      ,
    others => c_mgt_nil
    );

  constant c_REFCLK_TYPES : refclk_types_array_t (c_NUM_REFCLKS-1 downto 0) := (
    0      => REFCLK_SYNC320 ,
    1      => REFCLK_SYNC320 ,
    2      => REFCLK_SYNC320 ,
    3      => REFCLK_SYNC320 ,
    4      => REFCLK_SYNC320 ,
    others => REFCLK_NIL
    );

  -- FIXME: derive this constant in some sane way
  -- just make it oversized for now and the functions will just ignore the
  -- higher null values... make sure to only specify real things
  constant c_TDC_LINK_MAP : tdc_link_map_array_t (99*14-1 downto 0) := (
    -- TODO: we know that based on the CSM design (once it is final) there are
    -- only certain allowed pairs of even and odd elinks and these can be
    -- derived automatically by just specifying a slot number or something
    --
    -- this is assigned by the global MGT link ID (e.g. 0 to 75 on a ku15p)
    -- mgt link id           , even elink #, odd elink #, station
    0      => (link_id => 0   , even_elink => 0,  odd_elink => 1,  station_id => 0, legacy => false),
    1      => (link_id => 0   , even_elink => 2,  odd_elink => 3,  station_id => 0, legacy => false),
    2      => (link_id => 0   , even_elink => 4,  odd_elink => 5,  station_id => 0, legacy => false),
    3      => (link_id => 0   , even_elink => 6,  odd_elink => 7,  station_id => 0, legacy => false),
    4      => (link_id => 0   , even_elink => 8,  odd_elink => 9,  station_id => 0, legacy => false),
    5      => (link_id => 0   , even_elink => 10, odd_elink => 11, station_id => 0, legacy => false),
    6      => (link_id => 0   , even_elink => 12, odd_elink => 13, station_id => 0, legacy => false),
    7      => (link_id => 0   , even_elink => 14, odd_elink => 15, station_id => 0, legacy => false),
    8      => (link_id => 0   , even_elink => 16, odd_elink => 17, station_id => 0, legacy => false),
    9      => (link_id => 0   , even_elink => 18, odd_elink => 19, station_id => 0, legacy => false),
    10     => (link_id => 0   , even_elink => 20, odd_elink => 21, station_id => 0, legacy => false),
    11     => (link_id => 0   , even_elink => 22, odd_elink => 23, station_id => 0, legacy => false),
    12     => (link_id => 0   , even_elink => 24, odd_elink => 25, station_id => 0, legacy => false),
    13     => (link_id => 0   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    14     => (link_id => 1   , even_elink => 0,  odd_elink => 1,  station_id => 0, legacy => false),
    15     => (link_id => 1   , even_elink => 2,  odd_elink => 3,  station_id => 0, legacy => false),
    16     => (link_id => 1   , even_elink => 4,  odd_elink => 5,  station_id => 0, legacy => false),
    17     => (link_id => 1   , even_elink => 6,  odd_elink => 7,  station_id => 0, legacy => false),
    18     => (link_id => 1   , even_elink => 8,  odd_elink => 9,  station_id => 0, legacy => false),
    19     => (link_id => 1   , even_elink => 10, odd_elink => 11, station_id => 0, legacy => false),
    20     => (link_id => 1   , even_elink => 12, odd_elink => 13, station_id => 0, legacy => false),
    21     => (link_id => 1   , even_elink => 14, odd_elink => 15, station_id => 0, legacy => false),
    22     => (link_id => 1   , even_elink => 16, odd_elink => 17, station_id => 0, legacy => false),
    23     => (link_id => 1   , even_elink => 18, odd_elink => 19, station_id => 0, legacy => false),
    24     => (link_id => 1   , even_elink => 20, odd_elink => 21, station_id => 0, legacy => false),
    25     => (link_id => 1   , even_elink => 22, odd_elink => 23, station_id => 0, legacy => false),
    26     => (link_id => 1   , even_elink => 24, odd_elink => 25, station_id => 0, legacy => false),
    27     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    28     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    29     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    30     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    31     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    32     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    33     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    34     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    35     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    36     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    37     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    38     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    39     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    40     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    41     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    42     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    43     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    44     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    45     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    46     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    47     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    48     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    49     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    50     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    51     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    52     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    53     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    54     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    55     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    56     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    57     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    58     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    59     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    60     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    61     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    62     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    63     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    64     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    65     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    66     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    67     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    68     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    69     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    70     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    71     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    72     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    73     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    74     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    75     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    76     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    77     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    78     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    79     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    80     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    81     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    82     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    83     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    84     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    85     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    86     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    87     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    88     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    89     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    90     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    91     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    92     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    93     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    94     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    95     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    96     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    97     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    98     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    99     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    100     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    101     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    102     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    103     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    104     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    105     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    106     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    107     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    108     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    109     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    110     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    111     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    112     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    113     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    114     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    115     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    116     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    117     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    118     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    119     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    120     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    121     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    122     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    123     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    124     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    125     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    126     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    127     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    128     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    129     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    130     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    131     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    132     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    133     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    134     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    135     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    136     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    137     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    138     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    139     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    140     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    141     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    142     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    143     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    144     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    145     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    146     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    147     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    148     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    149     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    150     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    151     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    152     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    153     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    154     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    155     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    156     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    157     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    158     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    159     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    160     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    161     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    162     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    163     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    164     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    165     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    166     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    167     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    168     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    169     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    170     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    171     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    172     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    173     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    174     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    175     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    176     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    177     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    178     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    179     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    180     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    181     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    182     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    183     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    184     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    185     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    186     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    187     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    188     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    189     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    190     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    191     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    192     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    193     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    194     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    195     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    196     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    197     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    198     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    199     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    200     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    201     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    202     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    203     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    204     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    205     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    206     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    207     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    208     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    209     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    210     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    211     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    212     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    213     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    214     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    215     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    216     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    217     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    218     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    219     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    220     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    221     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    222     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    223     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    224     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    225     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    226     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    227     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    228     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    229     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    230     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    231     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    232     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    233     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    234     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    235     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    236     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    237     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    238     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    239     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    240     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    241     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    242     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    243     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    244     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    245     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    246     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    247     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    248     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    249     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    250     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    251     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    252     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    253     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    254     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    255     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    256     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    257     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    258     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    259     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    260     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    261     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    262     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    263     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    264     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    265     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    266     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    267     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    268     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    269     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    270     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    271     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    272     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    273     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    274     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    275     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    276     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    277     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    278     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    279     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    280     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    281     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    282     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    283     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    284     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    285     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    286     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    287     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    288     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    289     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    290     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    291     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    292     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    293     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    294     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    295     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    296     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    297     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    298     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    299     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    300     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    301     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    302     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    303     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    304     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    305     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    306     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    307     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    308     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    309     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    310     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    311     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    312     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    313     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    314     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    315     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    316     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    317     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    318     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    319     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    320     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    321     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    322     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    323     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    324     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    325     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    326     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    327     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    328     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    329     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    330     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    331     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    332     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    333     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    334     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    335     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    336     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    337     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    338     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    339     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    340     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    341     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    342     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    343     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    344     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    345     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    346     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    347     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    348     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    349     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    350     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    351     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    352     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    353     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    354     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    355     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    356     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    357     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    358     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    359     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    360     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    361     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    362     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    363     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    364     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    365     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    366     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    367     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    368     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    369     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    370     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    371     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    372     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    373     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    374     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    375     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    376     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    377     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    378     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    379     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    380     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    381     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    382     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    383     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    384     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    385     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    386     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    387     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    388     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    389     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    390     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    391     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    392     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    393     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    394     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    395     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    396     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    397     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    398     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    399     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    400     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    401     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    402     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    403     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    404     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    405     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    406     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    407     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    408     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    409     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    410     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    411     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    412     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    413     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    414     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    415     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    416     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    417     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    418     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    419     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    420     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    421     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    422     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    423     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    424     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    425     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    426     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    427     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    428     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    429     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    430     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    431     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    432     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    433     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    434     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    435     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    436     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    437     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    438     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    439     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    440     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    441     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    442     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    443     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    444     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    445     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    446     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),

    447     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    448     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    449     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    450     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    451     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    452     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    453     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    454     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    455     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    456     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    457     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    458     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    459     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    460     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    461     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    462     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    463     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    464     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    465     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    466     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    467     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    468     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    469     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    470     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    471     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    472     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    473     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    474     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    475     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    476     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    477     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    478     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    479     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    480     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    481     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    482     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    483     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    484     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    485     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    486     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    487     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    488     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    489     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    490     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    491     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    492     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    493     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    494     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    495     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    496     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    497     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    498     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    499     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    500     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    501     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    502     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    503     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    504     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    505     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    506     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    507     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    508     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    509     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    510     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    511     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    512     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    513     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    514     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    515     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    516     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    517     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    518     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    519     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    520     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    521     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    522     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    523     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    524     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    525     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    526     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    527     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    528     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    529     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    530     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    531     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    532     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    533     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    534     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    535     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    536     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    537     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    538     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    539     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    540     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    541     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    542     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    543     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    544     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    545     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    546     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    547     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    548     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    549     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    550     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    551     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    552     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    553     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    554     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    555     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    556     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    557     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    558     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    559     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    560     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    561     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    562     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    563     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    564     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    565     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    566     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    567     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    568     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    569     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    570     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    571     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    572     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    573     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    574     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    575     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    576     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    577     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    578     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    579     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    580     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    581     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    582     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    583     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    584     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    585     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    586     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    587     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    588     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    589     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    590     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    591     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    592     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    593     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    594     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    595     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    596     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    597     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    598     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    599     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    600     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    601     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    602     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    603     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    604     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    605     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    606     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    607     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    608     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    609     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    610     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    611     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    612     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    613     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    614     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    615     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    616     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    617     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    618     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    619     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    620     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    621     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    622     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    623     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    624     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    625     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    626     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    627     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    628     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    629     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    630     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    631     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    632     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    633     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    634     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    635     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    636     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    637     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    638     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    639     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    640     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    641     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    642     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    643     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    644     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    645     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    646     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    647     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    648     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    649     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    650     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    651     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    652     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    653     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    654     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    655     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    656     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    657     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    658     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    659     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    660     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    661     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    662     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    663     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    664     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    665     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    666     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    667     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    668     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    669     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    670     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => false),
    others => (-1, -1, -1, -1, false)
    );

end package board_pkg;
