library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.board_pkg_common.all;

package board_pkg is

  constant c_NUM_MGTS                 : integer := 44 + 32;
  constant c_NUM_REFCLKS              : integer := (c_NUM_MGTS/4);

  constant c_MGT_MAP : mgt_inst_array_t (c_NUM_MGTS-1 downto 0) := (

-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    0      => (MGT_LPGBT         , 0      , GTH     , 0 , 0)  ,
    1      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 1)  ,
    2      => (MGT_LPGBT         , 0      , GTH     , 0 , 2)  ,
    3      => (MGT_LPGBT_SIMPLEX , 0      , GTH     , 0 , 3)  ,
    4      => (MGT_LPGBT         , 1      , GTH     , 0 , 4)  ,
    5      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 5)  ,
    6      => (MGT_LPGBT         , 1      , GTH     , 0 , 6)  ,
    7      => (MGT_LPGBT_SIMPLEX , 1      , GTH     , 0 , 7)  ,
    8      => (MGT_LPGBT         , 2      , GTH     , 0 , 8)  ,
    9      => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 9)  ,
    10     => (MGT_LPGBT         , 2      , GTH     , 0 , 10) ,
    11     => (MGT_LPGBT_SIMPLEX , 2      , GTH     , 0 , 11) ,
    12     => (MGT_LPGBT         , 3      , GTH     , 0 , 12) ,
    13     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 13) ,
    14     => (MGT_LPGBT         , 3      , GTH     , 0 , 14) ,
    15     => (MGT_LPGBT_SIMPLEX , 3      , GTH     , 0 , 15) ,
    16     => (MGT_LPGBT         , 4      , GTH     , 0 , 16) ,
    17     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 17) ,
    18     => (MGT_LPGBT         , 4      , GTH     , 0 , 18) ,
    19     => (MGT_LPGBT_SIMPLEX , 4      , GTH     , 0 , 19) ,
    20     => (MGT_LPGBT         , 5      , GTH     , 0 , 20) ,
    21     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 21) ,
    22     => (MGT_LPGBT         , 5      , GTH     , 0 , 22) ,
    23     => (MGT_LPGBT_SIMPLEX , 5      , GTH     , 0 , 23) ,
    24     => (MGT_LPGBT         , 6      , GTH     , 0 , 24) ,
    25     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 25) ,
    26     => (MGT_LPGBT         , 6      , GTH     , 0 , 26) ,
    27     => (MGT_LPGBT_SIMPLEX , 6      , GTH     , 0 , 27) ,
    28     => (MGT_LPGBT         , 7      , GTH     , 0 , 28) ,
    29     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 29) ,
    30     => (MGT_LPGBT         , 7      , GTH     , 0 , 30) ,
    31     => (MGT_LPGBT_SIMPLEX , 7      , GTH     , 0 , 31) ,
    32     => (MGT_SL            , 8      , GTH     , 0 , 32) ,
    33     => (MGT_SL            , 8      , GTH     , 0 , 33) ,
    34     => (MGT_SL            , 8      , GTH     , 0 , 34) ,
    35     => (MGT_SL            , 8      , GTH     , 0 , 35) ,
    36     => (MGT_SL            , 9      , GTH     , 0 , 36) ,
    37     => (MGT_SL            , 9      , GTH     , 0 , 37) ,
    38     => (MGT_SL            , 9      , GTH     , 0 , 38) ,
    39     => (MGT_SL            , 9      , GTH     , 0 , 39) ,
    40     => (MGT_SL            , 10     , GTH     , 0 , 40) ,
    41     => (MGT_SL            , 10     , GTH     , 0 , 41) ,
    42     => (MGT_SL            , 10     , GTH     , 0 , 42) ,
    43     => (MGT_SL            , 10     , GTH     , 0 , 43) ,
-- mgt#    => (mgt_type          , refclk , gt_type , x , y)
    44     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 0)  ,
    45     => (MGT_LPGBT         , 11     , GTY     , 0 , 1)  ,
    46     => (MGT_LPGBT_SIMPLEX , 11     , GTY     , 0 , 2)  ,
    47     => (MGT_LPGBT         , 11     , GTY     , 0 , 3)  ,
    48     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 4)  ,
    49     => (MGT_LPGBT         , 12     , GTY     , 0 , 5)  ,
    50     => (MGT_LPGBT_SIMPLEX , 12     , GTY     , 0 , 6)  ,
    51     => (MGT_LPGBT         , 12     , GTY     , 0 , 7)  ,
    52     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 8)  ,
    53     => (MGT_LPGBT         , 13     , GTY     , 0 , 9)  ,
    54     => (MGT_LPGBT_SIMPLEX , 13     , GTY     , 0 , 10) ,
    55     => (MGT_LPGBT         , 13     , GTY     , 0 , 11) ,
    56     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 12) ,
    57     => (MGT_LPGBT         , 14     , GTY     , 0 , 13) ,
    58     => (MGT_LPGBT_SIMPLEX , 14     , GTY     , 0 , 14) ,
    59     => (MGT_LPGBT         , 14     , GTY     , 0 , 15) ,
    60     => c_mgt_nil ,
    61     => c_mgt_nil ,
    62     => c_mgt_nil ,
    63     => c_mgt_nil ,
    64     => c_mgt_nil ,
    65     => c_mgt_nil ,
    66     => c_mgt_nil ,
    67     => c_mgt_nil ,
    68     => c_mgt_nil ,
    69     => c_mgt_nil ,
    70     => c_mgt_nil ,
    71     => c_mgt_nil ,
    72     => c_mgt_nil ,
    73     => c_mgt_nil ,
    74     => c_mgt_nil ,
    75     => c_mgt_nil      ,
    others => c_mgt_nil
    );

  constant c_REFCLK_TYPES : refclk_types_array_t (c_NUM_REFCLKS-1 downto 0) := (
    0      => REFCLK_SYNC320 ,
    1      => REFCLK_SYNC320 ,
    2      => REFCLK_SYNC320 ,
    3      => REFCLK_SYNC320 ,
    4      => REFCLK_SYNC320 ,
    others => REFCLK_NIL
    );

  -- FIXME: derive this constant in some sane way
  -- just make it oversized for now and the functions will just ignore the
  -- higher null values... make sure to only specify real things
  constant c_TDC_LINK_MAP : tdc_link_map_array_t (99*14-1 downto 0) := (
    -- TODO: we know that based on the CSM design (once it is final) there are
    -- only certain allowed pairs of even and odd elinks and these can be
    -- derived automatically by just specifying a slot number or something
    --
    -- this is assigned by the global MGT link ID (e.g. 0 to 75 on a ku15p)
    -- mgt link id           , even elink #, odd elink #, station
    0      => (link_id => 0   , even_elink => 0,  odd_elink => 1,  station_id => 0, legacy => true),
    1      => (link_id => 0   , even_elink => 2,  odd_elink => 3,  station_id => 0, legacy => true),
    2      => (link_id => 0   , even_elink => 4,  odd_elink => 5,  station_id => 0, legacy => true),
    3      => (link_id => 0   , even_elink => 6,  odd_elink => 7,  station_id => 0, legacy => true),
    4      => (link_id => 0   , even_elink => 8,  odd_elink => 9,  station_id => 0, legacy => true),
    5      => (link_id => 0   , even_elink => 10, odd_elink => 11, station_id => 0, legacy => true),
    6      => (link_id => 0   , even_elink => 12, odd_elink => 13, station_id => 0, legacy => true),
    7      => (link_id => 0   , even_elink => 14, odd_elink => 15, station_id => 0, legacy => true),
    8      => (link_id => 0   , even_elink => 16, odd_elink => 17, station_id => 0, legacy => true),
    9      => (link_id => 0   , even_elink => 18, odd_elink => 19, station_id => 0, legacy => true),
    10     => (link_id => 0   , even_elink => 20, odd_elink => 21, station_id => 0, legacy => true),
    11     => (link_id => 0   , even_elink => 22, odd_elink => 23, station_id => 0, legacy => true),
    12     => (link_id => 0   , even_elink => 24, odd_elink => 25, station_id => 0, legacy => true),
    13     => (link_id => 0   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    14     => (link_id => 1   , even_elink => 0,  odd_elink => 1,  station_id => 0, legacy => true),
    15     => (link_id => 1   , even_elink => 2,  odd_elink => 3,  station_id => 0, legacy => true),
    16     => (link_id => 1   , even_elink => 4,  odd_elink => 5,  station_id => 0, legacy => true),
    17     => (link_id => 1   , even_elink => 6,  odd_elink => 7,  station_id => 0, legacy => true),
    18     => (link_id => 1   , even_elink => 8,  odd_elink => 9,  station_id => 0, legacy => true),
    19     => (link_id => 1   , even_elink => 10, odd_elink => 11, station_id => 0, legacy => true),
    20     => (link_id => 1   , even_elink => 12, odd_elink => 13, station_id => 0, legacy => true),
    21     => (link_id => 1   , even_elink => 14, odd_elink => 15, station_id => 0, legacy => true),
    22     => (link_id => 1   , even_elink => 16, odd_elink => 17, station_id => 0, legacy => true),
    23     => (link_id => 1   , even_elink => 18, odd_elink => 19, station_id => 0, legacy => true),
    24     => (link_id => 1   , even_elink => 20, odd_elink => 21, station_id => 0, legacy => true),
    25     => (link_id => 1   , even_elink => 22, odd_elink => 23, station_id => 0, legacy => true),
    26     => (link_id => 1   , even_elink => 24, odd_elink => 25, station_id => 0, legacy => true),
    27     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    28     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    29     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    30     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    31     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    32     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    33     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    34     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    35     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    36     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    37     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    38     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    39     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    40     => (link_id => 2   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    41     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    42     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    43     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    44     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    45     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    46     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    47     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    48     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    49     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    50     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    51     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    52     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    53     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    54     => (link_id => 3   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    55     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    56     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    57     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    58     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    59     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    60     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    61     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    62     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    63     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    64     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    65     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    66     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    67     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    68     => (link_id => 4   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    69     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    70     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    71     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    72     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    73     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    74     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    75     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    76     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    77     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    78     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    79     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    80     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    81     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    82     => (link_id => 5   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    83     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    84     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    85     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    86     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    87     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    88     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    89     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    90     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    91     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    92     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    93     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    94     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    95     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    96     => (link_id => 6   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    97     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    98     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    99     => (link_id => 7   , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    100     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    101     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    102     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    103     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    104     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    105     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    106     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    107     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    108     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    109     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    110     => (link_id => 7  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    111     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    112     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    113     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    114     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    115     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    116     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    117     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    118     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    119     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    120     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    121     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    122     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    123     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    124     => (link_id => 8  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    125     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    126     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    127     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    128     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    129     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    130     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    131     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    132     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    133     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    134     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    135     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    136     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    137     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    138     => (link_id => 9  , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    139     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    140     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    141     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    142     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    143     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    144     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    145     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    146     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    147     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    148     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    149     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    150     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    151     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    152     => (link_id => 10 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    153     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    154     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    155     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    156     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    157     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    158     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    159     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    160     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    161     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    162     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    163     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    164     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    165     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    166     => (link_id => 11 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    167     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    168     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    169     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    170     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    171     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    172     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    173     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    174     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    175     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    176     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    177     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    178     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    179     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    180     => (link_id => 12 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    181     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    182     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    183     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    184     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    185     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    186     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    187     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    188     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    189     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    190     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    191     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    192     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    193     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    194     => (link_id => 13 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    195     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    196     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    197     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    198     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    199     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    200     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    201     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    202     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    203     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    204     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    205     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    206     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    207     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    208     => (link_id => 14 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    209     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    210     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    211     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    212     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    213     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    214     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    215     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    216     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    217     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    218     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    219     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    220     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    221     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    222     => (link_id => 15 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    223     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    224     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    225     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    226     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    227     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    228     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    229     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    230     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    231     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    232     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    233     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    234     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    235     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    236     => (link_id => 16 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    237     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    238     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    239     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    240     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    241     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    242     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    243     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    244     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    245     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    246     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    247     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    248     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    249     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    250     => (link_id => 17 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    251     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    252     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    253     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    254     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    255     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    256     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    257     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    258     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    259     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    260     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    261     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    262     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    263     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    264     => (link_id => 18 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    265     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    266     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    267     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    268     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    269     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    270     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    271     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    272     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    273     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    274     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    275     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    276     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    277     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    278     => (link_id => 19 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    279     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    280     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    281     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    282     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    283     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    284     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    285     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    286     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    287     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    288     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    289     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    290     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    291     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    292     => (link_id => 20 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    293     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    294     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    295     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    296     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    297     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    298     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    299     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    300     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    301     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    302     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    303     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    304     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    305     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    306     => (link_id => 21 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    307     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    308     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    309     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    310     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    311     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    312     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    313     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    314     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    315     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    316     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    317     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    318     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    319     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    320     => (link_id => 22 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    321     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    322     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    323     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    324     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    325     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    326     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    327     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    328     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    329     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    330     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    331     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    332     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    333     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    334     => (link_id => 23 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    335     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    336     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    337     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    338     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    339     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    340     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    341     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    342     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    343     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    344     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    345     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    346     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    347     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    348     => (link_id => 24 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    349     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    350     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    351     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    352     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    353     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    354     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    355     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    356     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    357     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    358     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    359     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    360     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    361     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    362     => (link_id => 25 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    363     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    364     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    365     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    366     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    367     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    368     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    369     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    370     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    371     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    372     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    373     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    374     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    375     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    376     => (link_id => 26 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    377     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    378     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    379     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    380     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    381     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    382     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    383     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    384     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    385     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    386     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    387     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    388     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    389     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    390     => (link_id => 27 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    391     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    392     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    393     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    394     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    395     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    396     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    397     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    398     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    399     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    400     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    401     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    402     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    403     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    404     => (link_id => 28 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    405     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    406     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    407     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    408     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    409     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    410     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    411     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    412     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    413     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    414     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    415     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    416     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    417     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    418     => (link_id => 29 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    419     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    420     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    421     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    422     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    423     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    424     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    425     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    426     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    427     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    428     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    429     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    430     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    431     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    432     => (link_id => 30 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    433     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    434     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    435     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    436     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    437     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    438     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    439     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    440     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    441     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    442     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    443     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    444     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    445     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    446     => (link_id => 31 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),

    447     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    448     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    449     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    450     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    451     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    452     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    453     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    454     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    455     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    456     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    457     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    458     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    459     => (link_id => 44 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    460     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    461     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    462     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    463     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    464     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    465     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    466     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    467     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    468     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    469     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    470     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    471     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    472     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    473     => (link_id => 45 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    474     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    475     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    476     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    477     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    478     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    479     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    480     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    481     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    482     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    483     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    484     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    485     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    486     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    487     => (link_id => 46 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    488     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    489     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    490     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    491     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    492     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    493     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    494     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    495     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    496     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    497     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    498     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    499     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    500     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    501     => (link_id => 47 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    502     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    503     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    504     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    505     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    506     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    507     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    508     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    509     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    510     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    511     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    512     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    513     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    514     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    515     => (link_id => 48 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    516     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    517     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    518     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    519     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    520     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    521     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    522     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    523     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    524     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    525     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    526     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    527     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    528     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    529     => (link_id => 49 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    530     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    531     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    532     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    533     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    534     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    535     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    536     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    537     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    538     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    539     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    540     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    541     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    542     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    543     => (link_id => 50 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    544     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    545     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    546     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    547     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    548     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    549     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    550     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    551     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    552     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    553     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    554     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    555     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    556     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    557     => (link_id => 51 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    558     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    559     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    560     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    561     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    562     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    563     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    564     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    565     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    566     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    567     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    568     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    569     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    570     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    571     => (link_id => 52 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    572     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    573     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    574     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    575     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    576     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    577     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    578     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    579     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    580     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    581     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    582     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    583     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    584     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    585     => (link_id => 53 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    586     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    587     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    588     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    589     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    590     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    591     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    592     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    593     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    594     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    595     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    596     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    597     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    598     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    599     => (link_id => 54 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    600     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    601     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    602     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    603     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    604     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    605     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    606     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    607     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    608     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    609     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    610     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    611     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    612     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    613     => (link_id => 55 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    614     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    615     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    616     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    617     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    618     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    619     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    620     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    621     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    622     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    623     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    624     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    625     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    626     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    627     => (link_id => 56 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    628     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    629     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    630     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    631     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    632     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    633     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    634     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    635     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    636     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    637     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    638     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    639     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    640     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    641     => (link_id => 57 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    642     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    643     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    644     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    645     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    646     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    647     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    648     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    649     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    650     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    651     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    652     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    653     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    654     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    655     => (link_id => 58 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    656     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    657     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    658     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    659     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    660     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    661     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    662     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    663     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    664     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    665     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    666     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    667     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    668     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    669     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    670     => (link_id => 59 , even_elink => 26, odd_elink => 27, station_id => 0, legacy => true),
    others => (-1, -1, -1, -1, false)
    );

end package board_pkg;
