--------------------------------------------------------------------------------
--  UMass , Physics Department
--  Guillermo Loustau de Linares
--  gloustau@cern.ch
--------------------------------------------------------------------------------  
--  Project: ATLAS L0MDT Trigger 
--  Module: Hit Processor 
--          drift time - radius
--  Description:
--
--------------------------------------------------------------------------------
--  Revisions:
--      14/02/2019  0.1     File created
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library shared_lib;
use shared_lib.cfg_pkg.all;
use shared_lib.common_pkg.all;

library hp_lib;
use hp_lib.hp_pkg.all;

entity hp_calc_dt2r_small is
  generic(
    radius      : integer
  );
  port (
    clk                 : in std_logic;
    Reset_b             : in std_logic;
    glob_en             : in std_logic;

    i_drift_time        : in unsigned(HP_DRIFT_TIME_LEN -1 downto 0);
    i_data_valid        : in std_logic;
    o_tube_radius       : out unsigned(MDT_RADIUS_LEN -1 downto 0)
    -- o_data_valid        : out std_logic
  );
end entity hp_calc_dt2r_small;

architecture beh of hp_calc_dt2r_small is

begin


  DT2R : process(clk,Reset_b)

  begin
    if Reset_b = '0' then
      o_tube_radius <= (others => '0');
      -- o_data_valid <= '0';
    elsif rising_edge(clk) then
      -- o_data_valid <= i_data_valid;
      if(i_data_valid = '1') then
        -------------------------
        -- start of autogenerated code
        -------------------------
        
        if to_integer(i_drift_time) < 10 then
          o_tube_radius <= to_unsigned(1 ,MDT_RADIUS_LEN);
        elsif to_integer(i_drift_time) < 20 then
          o_tube_radius <= to_unsigned(2,MDT_RADIUS_LEN);
        end if;

        -------------------------
        -- end of autogenerated code
        -------------------------
      end if;

    end if ;
  end process;

end architecture beh;
