
find_max_bin find_max_bin_inst(
				  .ap_clk(clk),
				  .ap_rst(ap_rst),
				  .ap_start(results_ap_start),
				  .ap_done(results_ap_done),
				  .ap_idle(results_ap_idle),
				  .ap_ready(results_ap_ready),
				  .roi_seed_theta_V(roi_seed_theta),
				  .roi_seed_r_V(roi_seed_r[8]),	.max_bin_count_0_V(max_bin_count[0]),
.max_bin_r_0_V(max_bin_r[0]),
.max_bin_count_1_V(max_bin_count[1]),
.max_bin_r_1_V(max_bin_r[1]),
.max_bin_count_2_V(max_bin_count[2]),
.max_bin_r_2_V(max_bin_r[2]),
.max_bin_count_3_V(max_bin_count[3]),
.max_bin_r_3_V(max_bin_r[3]),
.max_bin_count_4_V(max_bin_count[4]),
.max_bin_r_4_V(max_bin_r[4]),
.max_bin_count_5_V(max_bin_count[5]),
.max_bin_r_5_V(max_bin_r[5]),
.max_bin_count_6_V(max_bin_count[6]),
.max_bin_r_6_V(max_bin_r[6]),
.max_bin_count_7_V(max_bin_count[7]),
.max_bin_r_7_V(max_bin_r[7]),
.max_bin_count_8_V(max_bin_count[8]),
.max_bin_r_8_V(max_bin_r[8]),
.max_bin_count_9_V(max_bin_count[9]),
.max_bin_r_9_V(max_bin_r[9]),
.max_bin_count_10_V(max_bin_count[10]),
.max_bin_r_10_V(max_bin_r[10]),
.max_bin_count_11_V(max_bin_count[11]),
.max_bin_r_11_V(max_bin_r[11]),
.max_bin_count_12_V(max_bin_count[12]),
.max_bin_r_12_V(max_bin_r[12]),
.max_bin_count_13_V(max_bin_count[13]),
.max_bin_r_13_V(max_bin_r[13]),
.max_bin_count_14_V(max_bin_count[14]),
.max_bin_r_14_V(max_bin_r[14]),
.max_bin_count_15_V(max_bin_count[15]),
.max_bin_r_15_V(max_bin_r[15]),
.max_bin_count_16_V(max_bin_count[16]),
.max_bin_r_16_V(max_bin_r[16]),
.max_bin_count_17_V(max_bin_count[17]),
.max_bin_r_17_V(max_bin_r[17]),
.max_bin_count_18_V(max_bin_count[18]),
.max_bin_r_18_V(max_bin_r[18]),
.max_bin_count_19_V(max_bin_count[19]),
.max_bin_r_19_V(max_bin_r[19]),
.max_bin_count_20_V(max_bin_count[20]),
.max_bin_r_20_V(max_bin_r[20]),
.max_bin_count_21_V(max_bin_count[21]),
.max_bin_r_21_V(max_bin_r[21]),
.max_bin_count_22_V(max_bin_count[22]),
.max_bin_r_22_V(max_bin_r[22]),
.max_bin_count_23_V(max_bin_count[23]),
.max_bin_r_23_V(max_bin_r[23]),
.max_bin_count_24_V(max_bin_count[24]),
.max_bin_r_24_V(max_bin_r[24]),
.max_bin_count_25_V(max_bin_count[25]),
.max_bin_r_25_V(max_bin_r[25]),
.max_bin_count_26_V(max_bin_count[26]),
.max_bin_r_26_V(max_bin_r[26]),
.max_bin_count_27_V(max_bin_count[27]),
.max_bin_r_27_V(max_bin_r[27]),
.max_bin_count_28_V(max_bin_count[28]),
.max_bin_r_28_V(max_bin_r[28]),
.max_bin_count_29_V(max_bin_count[29]),
.max_bin_r_29_V(max_bin_r[29]),
.max_bin_count_30_V(max_bin_count[30]),
.max_bin_r_30_V(max_bin_r[30]),
.max_bin_count_31_V(max_bin_count[31]),
.max_bin_r_31_V(max_bin_r[31]),
.max_bin_count_32_V(max_bin_count[32]),
.max_bin_r_32_V(max_bin_r[32]),
.max_bin_count_33_V(max_bin_count[33]),
.max_bin_r_33_V(max_bin_r[33]),
.max_bin_count_34_V(max_bin_count[34]),
.max_bin_r_34_V(max_bin_r[34]),
.max_bin_count_35_V(max_bin_count[35]),
.max_bin_r_35_V(max_bin_r[35]),
.max_bin_count_36_V(max_bin_count[36]),
.max_bin_r_36_V(max_bin_r[36]),
.max_bin_count_37_V(max_bin_count[37]),
.max_bin_r_37_V(max_bin_r[37]),
.max_bin_count_38_V(max_bin_count[38]),
.max_bin_r_38_V(max_bin_r[38]),
.max_bin_count_39_V(max_bin_count[39]),
.max_bin_r_39_V(max_bin_r[39]),
.max_bin_count_40_V(max_bin_count[40]),
.max_bin_r_40_V(max_bin_r[40]),
.max_bin_count_41_V(max_bin_count[41]),
.max_bin_r_41_V(max_bin_r[41]),
.max_bin_count_42_V(max_bin_count[42]),
.max_bin_r_42_V(max_bin_r[42]),
.max_bin_count_43_V(max_bin_count[43]),
.max_bin_r_43_V(max_bin_r[43]),
.max_bin_count_44_V(max_bin_count[44]),
.max_bin_r_44_V(max_bin_r[44]),
.max_bin_count_45_V(max_bin_count[45]),
.max_bin_r_45_V(max_bin_r[45]),
.max_bin_count_46_V(max_bin_count[46]),
.max_bin_r_46_V(max_bin_r[46]),
.max_bin_count_47_V(max_bin_count[47]),
.max_bin_r_47_V(max_bin_r[47]),
.max_bin_count_48_V(max_bin_count[48]),
.max_bin_r_48_V(max_bin_r[48]),
.max_bin_count_49_V(max_bin_count[49]),
.max_bin_r_49_V(max_bin_r[49]),
.max_bin_count_50_V(max_bin_count[50]),
.max_bin_r_50_V(max_bin_r[50]),
.max_bin_count_51_V(max_bin_count[51]),
.max_bin_r_51_V(max_bin_r[51]),
.max_bin_count_52_V(max_bin_count[52]),
.max_bin_r_52_V(max_bin_r[52]),
.max_bin_count_53_V(max_bin_count[53]),
.max_bin_r_53_V(max_bin_r[53]),
.max_bin_count_54_V(max_bin_count[54]),
.max_bin_r_54_V(max_bin_r[54]),
.max_bin_count_55_V(max_bin_count[55]),
.max_bin_r_55_V(max_bin_r[55]),
.max_bin_count_56_V(max_bin_count[56]),
.max_bin_r_56_V(max_bin_r[56]),
.max_bin_count_57_V(max_bin_count[57]),
.max_bin_r_57_V(max_bin_r[57]),
.max_bin_count_58_V(max_bin_count[58]),
.max_bin_r_58_V(max_bin_r[58]),
.max_bin_count_59_V(max_bin_count[59]),
.max_bin_r_59_V(max_bin_r[59]),
.max_bin_count_60_V(max_bin_count[60]),
.max_bin_r_60_V(max_bin_r[60]),
.max_bin_count_61_V(max_bin_count[61]),
.max_bin_r_61_V(max_bin_r[61]),
.max_bin_count_62_V(max_bin_count[62]),
.max_bin_r_62_V(max_bin_r[62]),
.max_bin_count_63_V(max_bin_count[63]),
.max_bin_r_63_V(max_bin_r[63]),
.max_bin_count_64_V(max_bin_count[64]),
.max_bin_r_64_V(max_bin_r[64]),
.max_bin_count_65_V(max_bin_count[65]),
.max_bin_r_65_V(max_bin_r[65]),
.max_bin_count_66_V(max_bin_count[66]),
.max_bin_r_66_V(max_bin_r[66]),
.max_bin_count_67_V(max_bin_count[67]),
.max_bin_r_67_V(max_bin_r[67]),
.max_bin_count_68_V(max_bin_count[68]),
.max_bin_r_68_V(max_bin_r[68]),
.max_bin_count_69_V(max_bin_count[69]),
.max_bin_r_69_V(max_bin_r[69]),
.max_bin_count_70_V(max_bin_count[70]),
.max_bin_r_70_V(max_bin_r[70]),
.max_bin_count_71_V(max_bin_count[71]),
.max_bin_r_71_V(max_bin_r[71]),
.max_bin_count_72_V(max_bin_count[72]),
.max_bin_r_72_V(max_bin_r[72]),
.max_bin_count_73_V(max_bin_count[73]),
.max_bin_r_73_V(max_bin_r[73]),
.max_bin_count_74_V(max_bin_count[74]),
.max_bin_r_74_V(max_bin_r[74]),
.max_bin_count_75_V(max_bin_count[75]),
.max_bin_r_75_V(max_bin_r[75]),
.max_bin_count_76_V(max_bin_count[76]),
.max_bin_r_76_V(max_bin_r[76]),
.max_bin_count_77_V(max_bin_count[77]),
.max_bin_r_77_V(max_bin_r[77]),
.max_bin_count_78_V(max_bin_count[78]),
.max_bin_r_78_V(max_bin_r[78]),
.max_bin_count_79_V(max_bin_count[79]),
.max_bin_r_79_V(max_bin_r[79]),
.max_bin_count_80_V(max_bin_count[80]),
.max_bin_r_80_V(max_bin_r[80]),
.max_bin_count_81_V(max_bin_count[81]),
.max_bin_r_81_V(max_bin_r[81]),
.max_bin_count_82_V(max_bin_count[82]),
.max_bin_r_82_V(max_bin_r[82]),
.max_bin_count_83_V(max_bin_count[83]),
.max_bin_r_83_V(max_bin_r[83]),
.max_bin_count_84_V(max_bin_count[84]),
.max_bin_r_84_V(max_bin_r[84]),
.max_bin_count_85_V(max_bin_count[85]),
.max_bin_r_85_V(max_bin_r[85]),
.max_bin_count_86_V(max_bin_count[86]),
.max_bin_r_86_V(max_bin_r[86]),
.max_bin_count_87_V(max_bin_count[87]),
.max_bin_r_87_V(max_bin_r[87]),
.max_bin_count_88_V(max_bin_count[88]),
.max_bin_r_88_V(max_bin_r[88]),
.max_bin_count_89_V(max_bin_count[89]),
.max_bin_r_89_V(max_bin_r[89]),
.max_bin_count_90_V(max_bin_count[90]),
.max_bin_r_90_V(max_bin_r[90]),
.max_bin_count_91_V(max_bin_count[91]),
.max_bin_r_91_V(max_bin_r[91]),
.max_bin_count_92_V(max_bin_count[92]),
.max_bin_r_92_V(max_bin_r[92]),
.max_bin_count_93_V(max_bin_count[93]),
.max_bin_r_93_V(max_bin_r[93]),
.max_bin_count_94_V(max_bin_count[94]),
.max_bin_r_94_V(max_bin_r[94]),
.max_bin_count_95_V(max_bin_count[95]),
.max_bin_r_95_V(max_bin_r[95]),
.max_bin_count_96_V(max_bin_count[96]),
.max_bin_r_96_V(max_bin_r[96]),
.max_bin_count_97_V(max_bin_count[97]),
.max_bin_r_97_V(max_bin_r[97]),
.max_bin_count_98_V(max_bin_count[98]),
.max_bin_r_98_V(max_bin_r[98]),
.max_bin_count_99_V(max_bin_count[99]),
.max_bin_r_99_V(max_bin_r[99]),
.max_bin_count_100_V(max_bin_count[100]),
.max_bin_r_100_V(max_bin_r[100]),
.max_bin_count_101_V(max_bin_count[101]),
.max_bin_r_101_V(max_bin_r[101]),
.max_bin_count_102_V(max_bin_count[102]),
.max_bin_r_102_V(max_bin_r[102]),
.max_bin_count_103_V(max_bin_count[103]),
.max_bin_r_103_V(max_bin_r[103]),
.max_bin_count_104_V(max_bin_count[104]),
.max_bin_r_104_V(max_bin_r[104]),
.max_bin_count_105_V(max_bin_count[105]),
.max_bin_r_105_V(max_bin_r[105]),
.max_bin_count_106_V(max_bin_count[106]),
.max_bin_r_106_V(max_bin_r[106]),
.max_bin_count_107_V(max_bin_count[107]),
.max_bin_r_107_V(max_bin_r[107]),
.max_bin_count_108_V(max_bin_count[108]),
.max_bin_r_108_V(max_bin_r[108]),
.max_bin_count_109_V(max_bin_count[109]),
.max_bin_r_109_V(max_bin_r[109]),
.max_bin_count_110_V(max_bin_count[110]),
.max_bin_r_110_V(max_bin_r[110]),
.max_bin_count_111_V(max_bin_count[111]),
.max_bin_r_111_V(max_bin_r[111]),
.max_bin_count_112_V(max_bin_count[112]),
.max_bin_r_112_V(max_bin_r[112]),
.max_bin_count_113_V(max_bin_count[113]),
.max_bin_r_113_V(max_bin_r[113]),
.max_bin_count_114_V(max_bin_count[114]),
.max_bin_r_114_V(max_bin_r[114]),
.max_bin_count_115_V(max_bin_count[115]),
.max_bin_r_115_V(max_bin_r[115]),
.max_bin_count_116_V(max_bin_count[116]),
.max_bin_r_116_V(max_bin_r[116]),
.max_bin_count_117_V(max_bin_count[117]),
.max_bin_r_117_V(max_bin_r[117]),
.max_bin_count_118_V(max_bin_count[118]),
.max_bin_r_118_V(max_bin_r[118]),
.max_bin_count_119_V(max_bin_count[119]),
.max_bin_r_119_V(max_bin_r[119]),
.max_bin_count_120_V(max_bin_count[120]),
.max_bin_r_120_V(max_bin_r[120]),
.max_bin_count_121_V(max_bin_count[121]),
.max_bin_r_121_V(max_bin_r[121]),
.max_bin_count_122_V(max_bin_count[122]),
.max_bin_r_122_V(max_bin_r[122]),
.max_bin_count_123_V(max_bin_count[123]),
.max_bin_r_123_V(max_bin_r[123]),
.max_bin_count_124_V(max_bin_count[124]),
.max_bin_r_124_V(max_bin_r[124]),
.max_bin_count_125_V(max_bin_count[125]),
.max_bin_r_125_V(max_bin_r[125]),
.max_bin_count_126_V(max_bin_count[126]),
.max_bin_r_126_V(max_bin_r[126]),
.max_bin_count_127_V(max_bin_count[127]),
.max_bin_r_127_V(max_bin_r[127]),
			       	  .hls_LT_theta_global_V(theta_global),
				  .hls_LT_theta_global_V_ap_vld(theta_global_vld),
				  .hls_LT_r_global_V(r_global),
				  .hls_LT_r_global_V_ap_vld(r_global_vld),
				  .hls_LT_theta_V(theta),
				  .hls_LT_theta_V_ap_vld(theta_vld),
				  .hls_LT_r_V(r),
				  .hls_LT_r_V_ap_vld(r_vld),
				  .res_max_bin_count_V(res_max_bin_count),
				  .res_max_bin_count_V_ap_vld(res_max_bin_count_vld),
				  .res_max_bin_theta_V(res_max_bin_theta),
				  .res_max_bin_theta_V_ap_vld(rest_max_bin_theta_vld),
				  .res_max_bin_r_V(res_max_bin_r),
				  .res_max_bin_r_V_ap_vld(res_max_bin_r_vld)
				  );
